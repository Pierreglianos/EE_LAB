library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;

package STATIC_MENU_PCKG is 
constant TECH_H_X_size : integer := 37;
constant TECH_H_Y_size : integer := 55;
type TECH_H_color_array is array(0 to TECH_H_Y_size - 1 , 0 to TECH_H_X_size - 1) of std_logic_vector(7 downto 0);

constant TECH_H_colors: TECH_H_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"6D", x"6D", x"49", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"DB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"6D", x"20"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"48", x"B6", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"48", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"48", x"49", x"6D", x"B6", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"91", x"B6", x"B6", x"BA", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"B6", x"B6", x"DA", x"DA", x"DB", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"DA", x"FF", x"FF", x"FF", x"FF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"20", x"48", x"DA", x"FF", x"FF", x"FF", x"FF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"24", x"24", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"24", x"49", x"6D", x"6D", x"91", x"DB", x"FF", x"FF", x"FF", x"FF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"6D", x"FF", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"24", x"71", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"24", x"71", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"24", x"71", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"24", x"91", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"24", x"91", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"24", x"91", x"DF", x"FF", x"FF", x"FF", x"DF", x"FF", x"FF", x"FF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"DF", x"FF", x"FF", x"DF", x"DF", x"FF", x"FF", x"6D", x"24"),
( x"24", x"91", x"DF", x"FF", x"DF", x"FF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"DF", x"FF", x"DF", x"FF", x"DF", x"DF", x"DF", x"FF", x"DF", x"6D", x"24"),
( x"24", x"91", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"B6", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"B6", x"91", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"91", x"B6", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BA", x"96", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"96", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"96", x"DF", x"DF", x"DF", x"DF", x"BF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"48", x"92", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"DF", x"BF", x"BF", x"BF", x"BF", x"BF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"DF", x"DF", x"DF", x"BF", x"DF", x"BF", x"DF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"DF", x"BF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"DF", x"BF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"72", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"72", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"72", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"71", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"6D", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"71", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"72", x"9F", x"9F", x"BF", x"9F", x"BF", x"9F", x"9F", x"9F", x"9F", x"6D", x"24"),
( x"24", x"6D", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"6D", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"72", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"6D", x"04"),
( x"00", x"49", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"72", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"48", x"00"),
( x"00", x"00", x"24", x"24", x"44", x"48", x"44", x"48", x"44", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"44", x"48", x"28", x"48", x"44", x"24", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);


constant FIGHTER_I_X_size : integer := 15;
constant FIGHTER_I_Y_size : integer := 54;
type FIGHTER_I_color_array is array(0 to FIGHTER_I_Y_size - 1 , 0 to FIGHTER_I_X_size - 1) of std_logic_vector(7 downto 0);

constant FIGHTER_I_colors: FIGHTER_I_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"B6", x"B6", x"B6", x"6E", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"DB", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"DB", x"FF", x"FF", x"FF", x"B7", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"DB", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00"),
( x"00", x"00", x"25", x"6D", x"6E", x"6E", x"92", x"DB", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00"),
( x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00"),
( x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6E", x"DF", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"FF", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6E", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6E", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6E", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"BB", x"DA", x"DB", x"DB", x"DB", x"D7", x"DB", x"DA", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B7", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"96", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"96", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"24", x"00", x"00"),
( x"00", x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"24", x"00", x"00"),
( x"00", x"04", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"24", x"00", x"00"),
( x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00"),
( x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"04", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"25", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

constant FIGHTER_H_X_size : integer := 36;
constant FIGHTER_H_Y_size : integer := 54;
type FIGHTER_H_color_array is array(0 to FIGHTER_H_Y_size - 1 , 0 to FIGHTER_H_X_size - 1) of std_logic_vector(7 downto 0);

constant FIGHTER_H_colors: FIGHTER_H_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6D", x"6D", x"6D", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"DB", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"DB", x"FF", x"FF", x"FF", x"DB", x"25"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"DB", x"FF", x"FF", x"FF", x"DB", x"25"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"49", x"49", x"DB", x"FF", x"FF", x"FF", x"DB", x"25"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6E", x"B6", x"B6", x"B7", x"B7", x"DB", x"FF", x"FF", x"FF", x"DB", x"25"),
( x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"DB", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"25"),
( x"00", x"00", x"00", x"00", x"00", x"49", x"DB", x"FF", x"FF", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"25"),
( x"00", x"00", x"00", x"00", x"25", x"6D", x"DB", x"FF", x"FF", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"25"),
( x"00", x"24", x"49", x"49", x"49", x"6E", x"DB", x"FF", x"FF", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"25"),
( x"00", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"DB", x"25"),
( x"24", x"B6", x"FF", x"DB", x"DF", x"FF", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"25"),
( x"24", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"25"),
( x"24", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"25"),
( x"24", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"BB", x"25"),
( x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"25"),
( x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"25"),
( x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"25"),
( x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25"),
( x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25"),
( x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25"),
( x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25"),
( x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25"),
( x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"6D", x"49", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"49", x"49", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25"),
( x"24", x"92", x"DA", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25"),
( x"24", x"92", x"DA", x"DB", x"B6", x"DB", x"DA", x"DB", x"BA", x"DA", x"DB", x"B6", x"DA", x"DA", x"B6", x"DA", x"BA", x"BA", x"DA", x"DA", x"BA", x"BA", x"DA", x"DA", x"B7", x"DB", x"DB", x"B7", x"DB", x"DB", x"B6", x"DB", x"DB", x"DB", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B7", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"BA", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"DB", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B7", x"B7", x"B7", x"B7", x"B7", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"6D", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"6D", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"96", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25"),
( x"24", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25"),
( x"24", x"92", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25"),
( x"24", x"92", x"92", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25"),
( x"24", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25"),
( x"24", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25"),
( x"24", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25"),
( x"24", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25"),
( x"24", x"8E", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"45"),
( x"24", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25"),
( x"24", x"6E", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6E", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25"),
( x"04", x"6E", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6E", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"24"),
( x"00", x"49", x"6D", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6D", x"24"),
( x"00", x"00", x"24", x"24", x"24", x"25", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00")
);


constant FIGHTER_T_X_size : integer := 40;
constant FIGHTER_T_Y_size : integer := 54;
type FIGHTER_T_color_array is array(0 to FIGHTER_T_Y_size - 1 , 0 to FIGHTER_T_X_size - 1) of std_logic_vector(7 downto 0);

constant FIGHTER_T_colors: FIGHTER_T_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"49"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"25", x"6E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49"),
( x"00", x"00", x"00", x"00", x"00", x"49", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6E", x"6E", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"DB", x"DB", x"B6", x"25"),
( x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"49", x"49", x"49", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"25", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"24", x"49", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"25", x"49", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"92", x"92", x"92", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"B6", x"B6", x"B6", x"B6", x"B2", x"B2", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00"),
( x"49", x"FF", x"FF", x"FF", x"DB", x"FF", x"DB", x"FF", x"DF", x"DB", x"DB", x"DB", x"FF", x"FF", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"25", x"24", x"24", x"24", x"24", x"24", x"24", x"20", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"69", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"6D", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"20", x"24", x"25", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B7", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B7", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"DA", x"B6", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"49", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

constant FIGHTER_F_X_size : integer := 34;
constant FIGHTER_F_Y_size : integer := 56;
type FIGHTER_F_color_array is array(0 to FIGHTER_F_Y_size - 1 , 0 to FIGHTER_F_X_size - 1) of std_logic_vector(7 downto 0);

constant FIGHTER_F_colors: FIGHTER_F_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"24", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6E", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"24", x"49", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"49", x"6D", x"6E", x"6E", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"DB", x"DB", x"92", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"69", x"49", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6E", x"25", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"04", x"25", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"25", x"49", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"6E", x"92", x"92", x"92", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"DB", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"DF", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"49", x"25", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"49", x"DB", x"DB", x"DB", x"FF", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DF", x"92", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"69", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"69", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"6E", x"6D", x"6D", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"69", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"69", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"69", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"69", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"69", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"49", x"24", x"20", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"DB", x"DA", x"D7", x"92", x"6E", x"6E", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"BB", x"DA", x"DB", x"DB", x"DB", x"D7", x"B6", x"B6", x"DB", x"B6", x"DB", x"DB", x"BA", x"DA", x"BA", x"DA", x"B6", x"DB", x"DB", x"DA", x"DA", x"B6", x"DA", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"D6", x"B7", x"BA", x"D7", x"B7", x"B6", x"B6", x"B6", x"DB", x"B6", x"BA", x"B6", x"B6", x"DB", x"B7", x"DB", x"B7", x"B6", x"B6", x"B7", x"B6", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B7", x"B7", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B7", x"B6", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"92", x"6E", x"25", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"49", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"6E", x"6E", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"96", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"92", x"B6", x"B2", x"92", x"96", x"B6", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"24", x"25", x"49", x"49", x"49", x"49", x"49", x"25", x"24", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

constant FIGHTER_G_X_size : integer := 37;
constant FIGHTER_G_Y_size : integer := 54;
type FIGHTER_G_color_array is array(0 to FIGHTER_G_Y_size - 1 , 0 to FIGHTER_G_X_size - 1) of std_logic_vector(7 downto 0);

constant FIGHTER_G_colors: FIGHTER_G_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"24", x"25", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"B6", x"B6", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"6E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"49", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"49", x"6E", x"6E", x"92", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"92", x"92", x"6E", x"49", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"49", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B7", x"DB", x"DB", x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"DB", x"92", x"92", x"92", x"92", x"B7", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"FF", x"FF", x"DB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"DB", x"FF", x"DB", x"FF", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"49", x"25", x"25", x"49", x"92", x"FF", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"FF", x"DB", x"B7", x"49", x"24", x"00", x"25", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00", x"00", x"00", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00", x"00", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"25", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"6D", x"6D", x"49", x"49", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"6D", x"6D", x"6D", x"6D", x"69", x"49", x"49", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"49", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"20", x"24", x"49", x"49", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"25", x"92", x"92", x"92", x"B2", x"B6", x"DA", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DA", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"B6", x"DB", x"DA", x"B7", x"DB", x"DB", x"DB", x"DA", x"B6", x"DB", x"B7", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"6D", x"BA", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"25", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"25", x"00", x"00"),
( x"00", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"6D", x"49", x"49", x"49", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"49", x"49", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"49", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6E", x"92", x"92", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00"),
( x"00", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"96", x"6D", x"25", x"24", x"00", x"00", x"00", x"00", x"24", x"25", x"6E", x"B6", x"B6", x"B2", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00"),
( x"24", x"6D", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"6E", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"6E", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"92", x"92", x"24", x"00"),
( x"24", x"69", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"96", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"49", x"49", x"25", x"00", x"00"),
( x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"49", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"25", x"49", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"49", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

constant FIGHTER_E_X_size : integer := 31;
constant FIGHTER_E_Y_size : integer := 54;
type FIGHTER_E_color_array is array(0 to FIGHTER_E_Y_size - 1 , 0 to FIGHTER_E_X_size - 1) of std_logic_vector(7 downto 0);

constant FIGHTER_E_colors: FIGHTER_E_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"24", x"25", x"24", x"24", x"24", x"04", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"B6", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B7", x"B6", x"B7", x"B6", x"B7", x"B6", x"92", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"6D", x"6E", x"6E", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"DB", x"B7", x"92", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"49", x"49", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"25", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6E", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"25", x"49", x"6E", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6E", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"6D", x"92", x"92", x"92", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"FF", x"DB", x"B6", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"B6", x"FF", x"DF", x"FF", x"DB", x"FF", x"DB", x"DB", x"DB", x"FB", x"DB", x"DB", x"FF", x"FF", x"B6", x"49", x"25", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"6D", x"49", x"49", x"45", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B7", x"49", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"25", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"DA", x"DB", x"DB", x"DA", x"DB", x"DB", x"DB", x"DB", x"B6", x"92", x"92", x"8E", x"8E", x"6E", x"6E", x"6E", x"8E", x"6E", x"8E", x"6E", x"6E", x"6E", x"6E", x"25", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"DA", x"DB", x"DB", x"DA", x"D7", x"DA", x"DA", x"DA", x"DB", x"B6", x"DB", x"B6", x"DA", x"DA", x"DA", x"BA", x"DA", x"DA", x"DA", x"DA", x"DB", x"B6", x"DB", x"6D", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B7", x"B6", x"B7", x"B6", x"B6", x"B7", x"B6", x"B6", x"BA", x"B6", x"D6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"20", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B7", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"20", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"8E", x"6E", x"6D", x"6D", x"25", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"6E", x"6D", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"45", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"25", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"45", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00"),
( x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"6D", x"24"),
( x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"96", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25"),
( x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49"),
( x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49"),
( x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"25"),
( x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"8E", x"6D", x"6D", x"49", x"49", x"20"),
( x"25", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"49", x"24", x"00", x"00", x"00"),
( x"25", x"6E", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"6D", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6E", x"6D", x"45", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

constant FIGHTER_R_X_size : integer := 32;
constant FIGHTER_R_Y_size : integer := 54;
type FIGHTER_R_color_array is array(0 to FIGHTER_R_Y_size - 1 , 0 to FIGHTER_R_X_size - 1) of std_logic_vector(7 downto 0);

constant FIGHTER_R_colors: FIGHTER_R_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"24", x"25", x"24", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"B6", x"B6", x"B7", x"B7", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"25", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B7", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B7", x"25", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B7", x"49", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6D", x"6D", x"6E", x"92", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"8E", x"6E", x"6D", x"49", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"49", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"00", x"00", x"24", x"25", x"49", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"25", x"92", x"92", x"92", x"92", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"B6", x"B6", x"B6", x"B7", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"49", x"FF", x"FF", x"DF", x"FB", x"DB", x"FF", x"DB", x"DB", x"DB", x"DB", x"FF", x"FF", x"DB", x"DB", x"6E", x"49", x"25", x"49", x"6E", x"DB", x"DB", x"FB", x"FF", x"DB", x"DB", x"DB", x"DB", x"FF", x"6D", x"00"),
( x"00", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"24", x"04", x"24", x"6E", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00", x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"04", x"6E", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"49", x"00", x"00", x"00", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"6E", x"6E", x"6D", x"49", x"24", x"00", x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6E", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6E", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6E", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"6E", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00"),
( x"24", x"6D", x"DA", x"DB", x"DB", x"DB", x"DB", x"DA", x"DA", x"DA", x"DA", x"6D", x"24", x"00", x"00", x"24", x"49", x"6D", x"6E", x"6E", x"92", x"B7", x"DB", x"DB", x"DB", x"DB", x"DA", x"DB", x"DA", x"DA", x"6D", x"04"),
( x"24", x"6D", x"B6", x"DB", x"DB", x"DB", x"D7", x"DA", x"DB", x"B7", x"B7", x"6D", x"00", x"00", x"00", x"49", x"B6", x"BA", x"BB", x"B7", x"B6", x"DB", x"BA", x"DA", x"DA", x"B6", x"DB", x"D7", x"B7", x"BB", x"6D", x"04"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B7", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"00", x"49", x"B6", x"B6", x"B6", x"DA", x"B6", x"B6", x"B6", x"DA", x"B6", x"DA", x"B6", x"B6", x"B6", x"BA", x"6D", x"04"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"24", x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B7", x"B7", x"B7", x"B6", x"B6", x"B7", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B7", x"B6", x"6E", x"49", x"25", x"49", x"6E", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"49", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"92", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"6E", x"6D", x"25", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"25", x"24", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"6D", x"6D", x"49", x"29", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"92", x"92", x"92", x"B6", x"B6", x"B6", x"B6", x"92", x"6E", x"6D", x"6D", x"49", x"25", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"49", x"49", x"49", x"6E", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6E", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"25", x"24", x"24", x"6D", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"25", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"24", x"00", x"24", x"49", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"49", x"24", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"6D", x"00", x"00", x"00", x"49", x"92", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"92", x"92", x"49", x"25", x"24", x"00", x"00", x"00"),
( x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"6E", x"6E", x"6D", x"25", x"00"),
( x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00"),
( x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00"),
( x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"04"),
( x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"04"),
( x"24", x"69", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"24", x"49", x"6D", x"6D", x"6E", x"8E", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00"),
( x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"45", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"24"),
( x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00"),
( x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00"),
( x"00", x"49", x"6D", x"6E", x"8E", x"92", x"8E", x"8E", x"92", x"6E", x"6D", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6D", x"6E", x"92", x"6E", x"92", x"92", x"8E", x"6E", x"6D", x"25", x"00"),
( x"00", x"00", x"24", x"25", x"25", x"25", x"25", x"25", x"25", x"25", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"25", x"25", x"25", x"25", x"25", x"25", x"24", x"24", x"00", x"00")
);

constant TECH_E_X_size : integer := 33;
constant TECH_E_Y_size : integer := 54;
type TECH_E_color_array is array(0 to TECH_E_Y_size - 1 , 0 to TECH_E_X_size - 1) of std_logic_vector(7 downto 0);

constant TECH_E_colors: TECH_E_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"20", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"48", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"44", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"91", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"28", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"48", x"4D", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"48", x"92", x"B6", x"B6", x"B6", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DA", x"B6", x"B6", x"6D", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"6D", x"48", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"96", x"48", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"48", x"91", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"6D", x"6D", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"71", x"20", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"96", x"92", x"91", x"91", x"91", x"91", x"91", x"91", x"6D", x"28", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"BA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"6D", x"48", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"48", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"48", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"DB", x"BA", x"BA", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"92", x"6D", x"48", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"DB", x"6D", x"24", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"FF", x"FF", x"FF", x"DF", x"DF", x"FF", x"FF", x"DB", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"FF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"6D", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"92", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"4D", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"DF", x"DF", x"DF", x"DB", x"DF", x"DF", x"DF", x"DB", x"DF", x"DF", x"DF", x"DF", x"DB", x"6D", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"BA", x"BB", x"BA", x"BA", x"6D", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"B6", x"6D", x"4D", x"48", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"B6", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"48", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"96", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"48", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"48", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"96", x"96", x"92", x"92", x"92", x"92", x"92", x"92", x"71", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"48", x"BA", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"6D", x"48", x"24", x"24", x"24", x"24", x"24", x"24", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"BF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BF", x"BB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"DF", x"BF", x"BB", x"49", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"DF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"6D", x"48", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00"),
( x"00", x"49", x"BA", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"B6", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"96", x"92", x"71", x"24", x"00"),
( x"00", x"49", x"9A", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00"),
( x"00", x"49", x"9A", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00"),
( x"00", x"49", x"9A", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00"),
( x"00", x"49", x"9A", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"9B", x"49", x"00"),
( x"00", x"49", x"9B", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"96", x"92", x"91", x"71", x"6D", x"24", x"00"),
( x"20", x"49", x"9A", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"96", x"49", x"24", x"24", x"00", x"00", x"00"),
( x"00", x"48", x"9A", x"9F", x"BF", x"BF", x"BF", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"92", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"28", x"7A", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"71", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"4D", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"76", x"49", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"04", x"24", x"24", x"28", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"48", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

constant TECH_C_X_size : integer := 37;
constant TECH_C_Y_size : integer := 55;
type TECH_C_color_array is array(0 to TECH_C_Y_size - 1 , 0 to TECH_C_X_size - 1) of std_logic_vector(7 downto 0);

constant TECH_C_colors: TECH_C_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"4D", x"4D", x"49", x"49", x"4D", x"49", x"6D", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"28", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"49", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"91", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"6D", x"48", x"24", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"92", x"B6", x"B6", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"B6", x"B6", x"92", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"48", x"49", x"6D", x"91", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"91", x"DB", x"DB", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"B6", x"92", x"92", x"92", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"91", x"48", x"48", x"49", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"6D", x"24", x"24", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"28", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"4D", x"20", x"00", x"24", x"91", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"24"),
( x"00", x"00", x"00", x"00", x"00", x"48", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"DF", x"DF", x"DF", x"DB", x"48", x"00", x"00", x"00", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"48", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"B6", x"6D", x"6D", x"49", x"48", x"24", x"00", x"00", x"00", x"24", x"48", x"49", x"6D", x"6D", x"6D", x"6D", x"6D", x"49", x"49", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"48", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"91", x"48", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"48", x"B6", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"48", x"B6", x"FF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"48", x"B6", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"48", x"B6", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"48", x"B6", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"49", x"B6", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"20", x"24", x"48", x"69", x"6D", x"B6", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"B6", x"BB", x"DB", x"DB", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"4D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"91", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"71", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"B6", x"6D", x"6D", x"49", x"44", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"96", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"48", x"72", x"92", x"96", x"96", x"96", x"96", x"96", x"92", x"71", x"24", x"00"),
( x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"BF", x"DF", x"DF", x"DF", x"6D", x"00"),
( x"24", x"6D", x"BF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"91", x"DF", x"DF", x"DF", x"DF", x"DF", x"BF", x"DF", x"BF", x"DF", x"6D", x"20"),
( x"24", x"6D", x"BF", x"BF", x"DF", x"BF", x"BF", x"DF", x"DF", x"BF", x"DF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"48", x"92", x"BF", x"BF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BF", x"6D", x"24"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"44", x"49", x"6D", x"96", x"DF", x"BF", x"BF", x"DF", x"BF", x"DF", x"DF", x"BF", x"DF", x"6D", x"24"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"BB", x"BB", x"BB", x"BB", x"BF", x"BF", x"BF", x"DF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"DF", x"BF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"24"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"96", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"48", x"91", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"6D", x"04"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"96", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"96", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"49", x"00"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BA", x"91", x"6D", x"69", x"49", x"24", x"00"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"9A", x"6D", x"44", x"24", x"00", x"00", x"00"),
( x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"96", x"48", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"4D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"96", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"96", x"9B", x"BB", x"9B", x"BB", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"9B", x"9A", x"9A", x"71", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"48", x"69", x"6D", x"96", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"9B", x"71", x"6D", x"48", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"49", x"96", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"9B", x"6D", x"24", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"96", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9B", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"52", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7B", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"28", x"4D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"49", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

constant TECH_T_X_size : integer := 42;
constant TECH_T_Y_size : integer := 55;
type TECH_T_color_array is array(0 to TECH_T_Y_size - 1 , 0 to TECH_T_X_size - 1) of std_logic_vector(7 downto 0);

constant TECH_T_colors: TECH_T_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"48", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"48", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"48", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"91", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"48", x"49", x"91", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"91", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"96", x"B6", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"DB", x"DB", x"B6", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"6D", x"49", x"24", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"48", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"48", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"6D", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"48", x"6D", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"B6", x"DB", x"DB", x"DB", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"96", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"48", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"4D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"6D", x"FF", x"DF", x"DF", x"DF", x"FF", x"FF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"91", x"92", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"48", x"71", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"FF", x"FF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"DF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"DF", x"BF", x"DF", x"DF", x"BF", x"BF", x"DF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"DF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"9B", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BB", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"BF", x"9B", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"9B", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9F", x"9A", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"7B", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"7F", x"76", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"4D", x"6D", x"71", x"71", x"71", x"71", x"71", x"6D", x"6D", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

constant TECH_Start_X 	: integer := 207;
constant TECH_End_X 		: integer := TECH_Start_X + TECH_T_X_size + TECH_E_X_size + TECH_C_X_size + TECH_H_X_size;
constant TECH_Start_Y 	: integer := 96;
constant TECH_End_Y 		: integer := TECH_Start_Y + TECH_H_Y_size;

constant FIGHTER_Start_X 	: integer := TECH_Start_X;
constant FIGHTER_End_X 		: integer := FIGHTER_Start_X + FIGHTER_F_X_size + FIGHTER_I_X_size + FIGHTER_G_X_size + FIGHTER_H_X_size + FIGHTER_T_X_size + FIGHTER_E_X_size + FIGHTER_R_X_size;
constant FIGHTER_Start_Y	: integer := TECH_End_Y + 30;
constant FIGHTER_End_Y		: integer := FIGHTER_Start_Y + FIGHTER_F_Y_size;

end STATIC_MENU_PCKG;