--library IEEE;
--use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--
--package player_renderer_package is
--
--constant PinkKick_X_size : integer := 44;
--constant PinkKick_Y_size : integer := 48;
--type PinkKick_color_array is array(0 to PinkKick_Y_size - 1 , 0 to PinkKick_X_size - 1) of std_logic_vector(7 downto 0);
--type PinkKick_bmp_array is array(0 to PinkKick_Y_size - 1 , 0 to PinkKick_X_size - 1) of std_logic;
--constant PinkKick_colors: PinkKick_color_array := (
--( x"DA", x"D6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DA", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"D2", x"AD", x"AD", x"AC", x"D2", x"FF", x"FF", x"FF", x"FF", x"D6", x"88", x"84", x"84", x"8C", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"88", x"88", x"A8", x"88", x"84", x"B1", x"FA", x"D6", x"AD", x"84", x"88", x"88", x"88", x"88", x"84", x"D6", x"FF", x"DB", x"B6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"88", x"88", x"88", x"88", x"88", x"88", x"A4", x"84", x"64", x"88", x"88", x"A8", x"A9", x"A9", x"A9", x"AD", x"D6", x"88", x"64", x"D1", x"D1", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"DA", x"B1", x"AD", x"DB", x"FB", x"FB", x"CD", x"A8", x"AC", x"A8", x"CD", x"AD", x"89", x"F6", x"F6", x"CD", x"A8", x"CD", x"AC", x"AD", x"AC", x"D1", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"F6", x"F2", x"F2", x"F2", x"89", x"8D", x"F6", x"FA", x"FA", x"FA", x"F1", x"AD", x"A8", x"CD", x"CD", x"CD", x"CC", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DB"),
--( x"DA", x"FF", x"FB", x"F2", x"F2", x"F7", x"F7", x"F7", x"F2", x"89", x"00", x"D5", x"F5", x"F5", x"F6", x"F6", x"F5", x"CD", x"88", x"64", x"B1", x"D6", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"D1"),
--( x"FF", x"FF", x"F2", x"ED", x"F2", x"F7", x"F7", x"F7", x"F2", x"89", x"00", x"D1", x"F5", x"F6", x"F6", x"F6", x"F6", x"F5", x"CD", x"8D", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F1", x"F6"),
--( x"FF", x"FB", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"CE", x"20", x"AD", x"F5", x"F6", x"FA", x"FA", x"F6", x"F5", x"F1", x"F5", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F5", x"F1"),
--( x"FF", x"F7", x"F7", x"EE", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"65", x"44", x"D1", x"F5", x"F6", x"F6", x"F5", x"FA", x"F6", x"F6", x"F5", x"F6", x"D2", x"69", x"64", x"89", x"8D", x"88", x"88", x"88", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"F5", x"F1", x"D1"),
--( x"FF", x"F6", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"D7", x"F2", x"CE", x"20", x"44", x"AD", x"F1", x"F6", x"F5", x"F5", x"F6", x"FA", x"FA", x"F5", x"64", x"40", x"40", x"40", x"40", x"40", x"40", x"60", x"CD", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F1", x"F5", x"F5", x"F1", x"D1"),
--( x"FF", x"F2", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"D2", x"69", x"64", x"AD", x"F5", x"F5", x"F5", x"F6", x"F6", x"F5", x"D1", x"60", x"60", x"40", x"40", x"60", x"40", x"40", x"60", x"F1", x"D1", x"FF", x"FF", x"FB", x"FB", x"FF", x"DA", x"D1", x"F1", x"F1", x"F5", x"F1", x"D1"),
--( x"FF", x"F2", x"F2", x"F7", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"F7", x"F2", x"EE", x"EE", x"C9", x"CD", x"ED", x"F1", x"F1", x"F1", x"D1", x"60", x"40", x"60", x"40", x"40", x"40", x"40", x"64", x"CD", x"D2", x"FB", x"F7", x"F7", x"F7", x"F7", x"F6", x"F1", x"F1", x"F1", x"F1", x"F5", x"F1"),
--( x"FF", x"F2", x"EE", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F2", x"EE", x"F2", x"EE", x"EE", x"C9", x"D1", x"D6", x"D6", x"FF", x"FF", x"B2", x"40", x"40", x"60", x"AD", x"AD", x"A8", x"CD", x"AC", x"D2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F5", x"F1", x"CD", x"F1", x"F1", x"CD"),
--( x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"AE", x"D2", x"F7", x"F7", x"D6", x"F6", x"D6", x"D7", x"F7", x"F7", x"F6", x"F7", x"F7", x"F2", x"F1", x"D2", x"D6", x"FA", x"FB", x"FB"),
--( x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F2", x"EE", x"CD", x"A9", x"89", x"C9", x"EE", x"FF", x"FF", x"FB", x"F7", x"F7", x"F7", x"FB", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F3", x"EE", x"A9", x"64", x"44", x"64", x"44", x"A9", x"EE", x"F2", x"F7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"69", x"20", x"40", x"89", x"AE", x"CE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"89", x"20", x"89", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B2", x"D2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"F2", x"EE", x"EE", x"F2", x"F6", x"F6", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F7", x"F7", x"D7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"EE", x"F2", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"C9", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F6", x"F2", x"EE", x"EE", x"E9", x"EE", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"F2", x"F2", x"F7", x"D7", x"F7", x"F2", x"EE", x"E9", x"C9", x"C9", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"EE", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"EE", x"ED", x"CD", x"ED", x"F2", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"CE", x"C9", x"CD", x"CD", x"ED", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F6", x"CD", x"F1", x"F1", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"CD", x"F5", x"F1", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F1", x"F5", x"F5", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F1", x"F1", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"CD", x"AD", x"AC", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"CD", x"F1", x"CD", x"CD", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CC", x"CD", x"CD", x"CD", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
--);
--constant PinkKick_bmp: PinkKick_bmp_array := (
--("11100000001110000000000000000000000000000000"),
--("11111000011111100000000000000000000000000000"),
--("11111111111111110111000000000000000000000000"),
--("11111111111111111111110000000000000000000000"),
--("11111111111111111111111100000000000000000000"),
--("01000011111111111111111100000000000000000011"),
--("10111111111111111111111100000000000000000111"),
--("00111111111111111111100000000000000000001111"),
--("01111111111111111111100000000000000000001111"),
--("01111111111111111111111111111110000000011111"),
--("01111111111111111111111111111111000000111111"),
--("01111111111111111111111111111111001101111111"),
--("01111111111111111111111111111111111111111111"),
--("01111111111111111111001111111111111111111111"),
--("00111111111111111100000111111111111111111111"),
--("00011111111111111001111111111111111111100000"),
--("00001111111111111111111111111111111111100000"),
--("00000111111111111111111111111111111000000000"),
--("00000011111111111111111111111111100000000000"),
--("00000011111111111111111111111110000000000000"),
--("00000011111111111111111110000000000000000000"),
--("00000011111111111111111100000000000000000000"),
--("00000011111111111111110000000000000000000000"),
--("00000011111111111111000000000000000000000000"),
--("00000001111111111100000000000000000000000000"),
--("00000001111111111000000000000000000000000000"),
--("00000001111111111000000000000000000000000000"),
--("00000001111111110000000000000000000000000000"),
--("00000001111111110000000000000000000000000000"),
--("00000001111111110000000000000000000000000000"),
--("00000001111111100000000000000000000000000000"),
--("00000001111111100000000000000000000000000000"),
--("00000011111111100000000000000000000000000000"),
--("00000011111111100000000000000000000000000000"),
--("00000011111111000000000000000000000000000000"),
--("00000011111111000000000000000000000000000000"),
--("00000011111111000000000000000000000000000000"),
--("00000011111111000000000000000000000000000000"),
--("00000011111110000000000000000000000000000000"),
--("00000111111110000000000000000000000000000000"),
--("00000111111100000000000000000000000000000000"),
--("00000011111100000000000000000000000000000000"),
--("00000001111100000000000000000000000000000000"),
--("00000001111100000000000000000000000000000000"),
--("00000001111100000000000000000000000000000000"),
--("00000011111100000000000000000000000000000000"),
--("00000111111100000000000000000000000000000000"),
--("00000111111100000000000000000000000000000000")
--);
--constant PinkDucking_X_size : integer := 53;
--constant PinkDucking_Y_size : integer := 48;
--type PinkDucking_color_array is array(0 to PinkDucking_Y_size - 1 , 0 to PinkDucking_X_size - 1) of std_logic_vector(7 downto 0);
--type PinkDucking_bmp_array is array(0 to PinkDucking_Y_size - 1 , 0 to PinkDucking_X_size - 1) of std_logic;
--constant PinkDucking_colors: PinkDucking_color_array := (
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"D1", x"B1", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"8D", x"84", x"84", x"88", x"88", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"88", x"88", x"A8", x"88", x"88", x"AC", x"AC", x"84", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"F7", x"D2", x"A8", x"88", x"AC", x"D1", x"D1", x"AD", x"44", x"F5", x"AC", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"F7", x"F2", x"F2", x"EE", x"EE", x"C9", x"C9", x"CD", x"ED", x"F1", x"CD", x"D5", x"FA", x"F6", x"AD", x"CD", x"D2", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"D2", x"D2", x"F2", x"F2", x"EE", x"F3", x"D2", x"CD", x"F1", x"F5", x"F1", x"F1", x"CD", x"F5", x"FA", x"F6", x"D1", x"D1", x"F2", x"D2", x"F7", x"F2", x"D2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F5", x"F6", x"F2", x"F7", x"F3", x"F2", x"F7", x"A9", x"68", x"F1", x"F5", x"F5", x"F1", x"F1", x"AC", x"D1", x"D1", x"CD", x"F2", x"F7", x"F7", x"F2", x"EE", x"CD", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F2", x"F2", x"F7", x"F3", x"F2", x"F7", x"A9", x"00", x"48", x"68", x"44", x"68", x"44", x"00", x"89", x"F2", x"EE", x"F7", x"D7", x"F7", x"F2", x"F1", x"FA", x"F1", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F1", x"F2", x"F7", x"F7", x"F2", x"F7", x"AD", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"89", x"F7", x"EE", x"F2", x"F7", x"F2", x"F1", x"F5", x"F5", x"D1", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F2", x"F2", x"F7", x"EE", x"F7", x"B2", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"D2", x"F3", x"F2", x"F7", x"F2", x"CD", x"F1", x"FA", x"F6", x"F5", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"EE", x"F2", x"F7", x"F2", x"F2", x"F7", x"65", x"00", x"00", x"20", x"45", x"8E", x"D2", x"F7", x"F2", x"F7", x"F7", x"EE", x"CD", x"CD", x"F5", x"FA", x"FA", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"D6", x"A8", x"A8", x"C9", x"C9", x"F2", x"F2", x"EE", x"F6", x"D7", x"69", x"44", x"D2", x"F3", x"F2", x"F2", x"EE", x"F6", x"F3", x"F2", x"F2", x"CD", x"AD", x"CD", x"D1", x"F6", x"F5", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FA", x"FB", x"FB", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"D1", x"CD", x"AC", x"AC", x"A8", x"CD", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"ED", x"CD", x"F1", x"CD", x"CD", x"CD", x"F1", x"D1", x"D1", x"F6", x"FA", x"FB", x"D6", x"D6", x"B6", x"D6", x"D6", x"F5", x"A8", x"8C", x"8D", x"D1", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"AD", x"D1", x"F1", x"F5", x"F1", x"CD", x"A9", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"ED", x"EE", x"F6", x"DA", x"B1", x"A8", x"D1", x"D1", x"F5", x"F6", x"F5", x"F5", x"F5", x"F5", x"D1", x"40", x"40", x"60", x"D1", x"D1", x"64", x"B1", x"D1", x"B1", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"8D", x"88", x"88", x"88", x"A8", x"64", x"20", x"44", x"A9", x"C9", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"C9", x"C9", x"CD", x"F6", x"FB", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"F5", x"F6", x"F6", x"F5", x"F5", x"F6", x"D1", x"40", x"40", x"40", x"D1", x"F1", x"68", x"D1", x"D1", x"DA", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D2", x"CE", x"CD", x"EE", x"85", x"40", x"20", x"20", x"60", x"65", x"65", x"64", x"60", x"64", x"40", x"A9", x"F2", x"FB", x"FB", x"F6", x"FB", x"FF", x"FF", x"D6", x"D6", x"F6", x"D6", x"D6", x"D6", x"D1", x"D1", x"AD", x"64", x"40", x"40", x"88", x"AC", x"44", x"64", x"AD", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"F7", x"F7", x"F7", x"F7", x"F3", x"F2", x"F2", x"EE", x"EE", x"CE", x"AD", x"65", x"00", x"00", x"00", x"89", x"C9", x"CD", x"F2", x"F2", x"EE", x"F7", x"F2", x"F7", x"F7", x"F7", x"FB", x"FF", x"FB", x"FB", x"F7", x"FB", x"FF", x"FF", x"FF", x"FB", x"D6", x"FB", x"DB", x"D6", x"D6", x"D6", x"DB", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FB", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"F2", x"CE", x"24", x"44", x"A9", x"20", x"69", x"EE", x"EE", x"EE", x"F2", x"D7", x"F7", x"F7", x"F7", x"F7", x"D7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F2", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"65", x"00", x"C9", x"EE", x"65", x"00", x"A9", x"EE", x"EE", x"F2", x"F6", x"F2", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"F2", x"F7", x"D7", x"F3", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"F6", x"EE", x"F2", x"F7", x"F2", x"F7", x"F6", x"F2", x"F2", x"EE", x"F2", x"F7", x"F2", x"EE", x"EE", x"EE", x"24", x"24", x"E9", x"EE", x"A9", x"00", x"85", x"EE", x"EE", x"EE", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"F7", x"F7", x"F7", x"F2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F7", x"F2", x"CE", x"C9", x"F2", x"F2", x"EE", x"EE", x"A9", x"00", x"85", x"E9", x"E9", x"E9", x"40", x"20", x"EA", x"EE", x"EE", x"EE", x"F2", x"EE", x"E9", x"EE", x"EE", x"EE", x"EE", x"F2", x"F7", x"F7", x"F6", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"EE", x"F2", x"EE", x"F2", x"EE", x"EE", x"F2", x"F7", x"EE", x"CE", x"EE", x"EE", x"F2", x"F2", x"AD", x"00", x"A9", x"D2", x"EE", x"F2", x"44", x"20", x"F2", x"F2", x"F2", x"F2", x"F2", x"D2", x"D2", x"F6", x"CE", x"C5", x"EE", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"96", x"DB", x"FF", x"FF", x"FF", x"B6", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F7", x"F2", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EA", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F3", x"F7", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"F2", x"CD", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"EE", x"EE", x"EE", x"EE", x"ED", x"CE", x"F7", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FB", x"D1", x"CD", x"F1", x"ED", x"ED", x"F2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F6", x"CD", x"CD", x"CD", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"F2", x"F1", x"F5", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"CD", x"F1", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FA", x"F5", x"F1", x"F1", x"F1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D6", x"F1", x"F1", x"F1", x"F5", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"F1", x"F5", x"F5", x"F1", x"F5", x"F1", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"D6", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"D1", x"F1", x"F5", x"F5", x"F1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"D1", x"F1", x"F1", x"F1", x"F1", x"F1", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F1", x"F5", x"F1", x"F1", x"D1", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"D5", x"F6", x"D6", x"F6", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FA", x"FB", x"FA", x"FA", x"FA", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
--);
--constant PinkDucking_bmp: PinkDucking_bmp_array := (
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000000000000000000"),
--("00000000000000000000000001111100000000000000000000000"),
--("00000000000000000000000111111110000000000000000000000"),
--("00000000000000000000001111111111000000000000000000000"),
--("00000000000000000011111111111111000000000000000000000"),
--("00000000000011111111111111111111000000000000000000000"),
--("00000000000111111111111111111111111100000000000000000"),
--("00000000001111111111111111111111111110000000000000000"),
--("00000000001111111111111111111111111110000000000000000"),
--("00000000000111111111111111111111111110000000000000000"),
--("00000000000111111111111111111111111110000000000000000"),
--("00000000000111111111111111111111111110000000000000000"),
--("00000000011111111111111111111111111111100000000111100"),
--("00000000111111111111111111111111111111111111111111110"),
--("00000000111111111111111111111111111111111111111111110"),
--("00000000011111111111111111111100011111111111111111110"),
--("00000000001111111111111111111111001111111111111111100"),
--("00000011111111111111111111111111111011110001111111100"),
--("00011111111111111111111111111111111111111100000000000"),
--("00111111111111111111111111111111111111111100000000000"),
--("00111111111111111111111111111111111111111100000000000"),
--("00111111111111111111111111111111111111111110000000000"),
--("00111111111111111111111111111111111111111110000000000"),
--("00111111111110000011000110000000011111111111000000000"),
--("00011111111100000000000000000000011111111111100000000"),
--("00011111111100000000000000000000001111111111100000000"),
--("00011111111000000000000000000000000111111100000000000"),
--("00001111100000000000000000000000000011111000000000000"),
--("00011111100000000000000000000000001111111000000000000"),
--("00111111110000000000000000000000001111111100000000000"),
--("01111111110000000000000000000000001111111100000000000"),
--("11111111000000000000000000000000000001111111110000000"),
--("11111100000000000000000000000000000000111111110000000")
--);
--constant PinkHitted_X_size : integer := 38;
--constant PinkHitted_Y_size : integer := 48;
--type PinkHitted_color_array is array(0 to PinkHitted_Y_size - 1 , 0 to PinkHitted_X_size - 1) of std_logic_vector(7 downto 0);
--type PinkHitted_bmp_array is array(0 to PinkHitted_Y_size - 1 , 0 to PinkHitted_X_size - 1) of std_logic;
--constant PinkHitted_colors: PinkHitted_color_array := (
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FB", x"B1", x"8C", x"AD", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"88", x"AC", x"88", x"88", x"84", x"84", x"AD", x"FF", x"FF", x"FF", x"FB", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"B1", x"88", x"B1", x"D1", x"CC", x"88", x"AC", x"84", x"B1", x"FF", x"DA", x"AD", x"AD", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"A8", x"AC", x"48", x"D5", x"D5", x"AC", x"F6", x"A8", x"A8", x"AD", x"A8", x"84", x"B1", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"DB", x"B2", x"B1", x"AD", x"89", x"F1", x"F6", x"D1", x"F1", x"F1", x"D1", x"A8", x"88", x"88", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"CD", x"D1", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FB", x"FB", x"FF", x"D2", x"CD", x"F5", x"F6", x"FA", x"F6", x"F1", x"F5", x"F5", x"CD", x"CD", x"CE", x"CE", x"F6", x"F2", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"FF", x"B6", x"AD", x"CD", x"D1", x"CD", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"F6", x"D1", x"F6", x"F6", x"F5", x"D1", x"F5", x"F5", x"F6", x"F1", x"CD", x"88", x"A9", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F5", x"68", x"24", x"88", x"CD", x"CD", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"CD", x"D1", x"D2", x"F6", x"F6", x"F2", x"F1", x"F5", x"D1", x"88", x"20", x"85", x"EE", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F1", x"44", x"00", x"44", x"88", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"F2", x"E9", x"EE", x"EE", x"F2", x"F3", x"F7", x"F3", x"F7", x"F2", x"F1", x"64", x"00", x"00", x"85", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"DB", x"88", x"CD", x"CD", x"AC", x"48", x"00", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"F2", x"AD", x"89", x"D2", x"F2", x"F2", x"F2", x"F7", x"F3", x"F3", x"F2", x"F7", x"F3", x"8D", x"24", x"00", x"C9", x"F2", x"F1", x"FA", x"FB", x"FA", x"AC", x"20", x"40", x"64", x"C8", x"A8", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"F7", x"EA", x"65", x"68", x"69", x"49", x"69", x"F2", x"F7", x"F7", x"D7", x"D7", x"F7", x"F7", x"F6", x"F7", x"D2", x"44", x"40", x"CE", x"EE", x"CC", x"CD", x"F5", x"D1", x"60", x"20", x"20", x"20", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"F2", x"89", x"B5", x"FA", x"FA", x"F6", x"D1", x"8D", x"AE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"44", x"A9", x"EE", x"CD", x"F1", x"F1", x"F1", x"CC", x"A8", x"88", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"CE", x"8D", x"F5", x"FA", x"FA", x"F5", x"F1", x"F6", x"D1", x"F2", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"F2", x"D2", x"CE", x"EE", x"EE", x"CD", x"CD", x"ED", x"F1", x"F1", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"D2", x"A9", x"F1", x"F1", x"F5", x"F5", x"F5", x"F6", x"FA", x"F5", x"CD", x"EE", x"F2", x"F3", x"F7", x"F7", x"F7", x"EE", x"F2", x"F2", x"E9", x"EE", x"C9", x"CD", x"CD", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"CE", x"CD", x"F1", x"F1", x"F6", x"FA", x"F6", x"F5", x"F1", x"CD", x"CD", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"A5", x"A9", x"84", x"A5", x"C8", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FA", x"F1", x"F5", x"F5", x"F1", x"F5", x"F6", x"F6", x"F6", x"F5", x"F1", x"D1", x"CD", x"A9", x"64", x"60", x"40", x"40", x"20", x"8D", x"F5", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FA", x"D1", x"F5", x"F5", x"D1", x"F6", x"FA", x"F6", x"F6", x"FA", x"F6", x"84", x"40", x"40", x"40", x"60", x"40", x"64", x"F5", x"F6", x"F5", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"A9", x"F1", x"D1", x"CD", x"F5", x"F6", x"FA", x"FA", x"F6", x"60", x"40", x"40", x"40", x"60", x"40", x"AD", x"F6", x"F5", x"F1", x"D1", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"C9", x"F1", x"F5", x"F1", x"F1", x"F5", x"F5", x"F5", x"64", x"40", x"40", x"40", x"40", x"64", x"D1", x"D5", x"F5", x"CD", x"D1", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D6", x"D1", x"D1", x"F1", x"F1", x"F1", x"CD", x"CD", x"A9", x"84", x"85", x"C9", x"A9", x"20", x"44", x"AD", x"CD", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"CD", x"CD", x"C9", x"EE", x"F3", x"F2", x"F2", x"F2", x"F2", x"EE", x"00", x"40", x"20", x"89", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"C9", x"EE", x"EE", x"EE", x"F2", x"F7", x"F7", x"F2", x"EE", x"EA", x"40", x"20", x"44", x"00", x"A9", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"C9", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"ED", x"EE", x"A9", x"00", x"64", x"44", x"00", x"A9", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"EE", x"EE", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"E9", x"40", x"20", x"89", x"00", x"00", x"D2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EA", x"EE", x"85", x"00", x"69", x"AE", x"69", x"D7", x"F3", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"F7", x"F7", x"F7", x"D7", x"F7", x"F2", x"E9", x"F2", x"A9", x"20", x"AE", x"FB", x"F7", x"D7", x"F7", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"C9", x"EE", x"F2", x"D2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"CE", x"EE", x"EE", x"F2", x"F7", x"F2", x"F7", x"D7", x"F7", x"D7", x"F7", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"EE", x"F2", x"FB", x"EE", x"F2", x"F7", x"F7", x"F2", x"F7", x"D7", x"F7", x"F7", x"F2", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"EE", x"F2", x"FF", x"F2", x"EE", x"F2", x"F7", x"F7", x"F6", x"F7", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"EA", x"F3", x"F7", x"F7", x"F7", x"D7", x"F7", x"EE", x"F6", x"FF", x"FF", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"CE", x"FB", x"FF", x"FF", x"FF", x"F2", x"C9", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"F6", x"C9", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"E9", x"EE", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"F7", x"EA", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"E9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"E9", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F7", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"ED", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"D1", x"ED", x"ED", x"ED", x"F6", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"ED", x"ED", x"CD", x"F2", x"EE", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"CD", x"CD", x"F1", x"F5", x"F1", x"F6", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"F1", x"CD", x"CD", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"F1", x"F5", x"F5", x"F1", x"FB", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"F5", x"F5", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"F5", x"F5", x"F5", x"D1", x"FB"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F1", x"F5", x"F1", x"F1", x"F1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"D1", x"F1", x"D1", x"CD", x"D6"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"F1", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"D1", x"CD", x"CD", x"D6", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D2", x"D6", x"D2", x"D6", x"D2", x"D6", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"D6", x"FB", x"FF", x"FF")
--);
--constant PinkHitted_bmp: PinkHitted_bmp_array := (
--("00000000000000000000000000000000000000"),
--("00000000000000000000000000000000000000"),
--("00011111100001000000000000000000000000"),
--("00111111110001100000000000000000000000"),
--("00111111111011110000000000000000000000"),
--("01111111111111110000000000000100000000"),
--("11111111111111110000000000011111000000"),
--("11011111111111111111000001011111100000"),
--("00001111111111111111000001111111110000"),
--("00001111111111111111100000111111110000"),
--("00001111111111111111100001111111100000"),
--("00111111111111111111111111111111000000"),
--("01111111111111111111111111111110000000"),
--("01111111111111111111111111111100000000"),
--("01111111111111111111111111111000000000"),
--("01111111111111111111111111110000000000"),
--("01111111111111111111111111000000000000"),
--("00011111111111111111111111000000000000"),
--("00001111111111111111111111100000000000"),
--("00000111111111111111111111100000000000"),
--("00000011111111111111111111100000000000"),
--("00000001111111111111111111110000000000"),
--("00000000011111111111111111110000000000"),
--("00000000001111111111111111110000000000"),
--("00000000001111111111111111111000000000"),
--("00000000001111111111111111111000000000"),
--("00000000001111111111111111111100000000"),
--("00000000000111111111111111111110000000"),
--("00000000000111111111111111111111000000"),
--("00000000001111111111111111111111100000"),
--("00000000000111111111111111111111100000"),
--("00000000000111111111101111111111100000"),
--("00000000001111111111100111111111110000"),
--("00000000001111111111100011111111110000"),
--("00000000001111111111100011111111110000"),
--("00000000011111111111000011111111110000"),
--("00000000011111111111000001111111111000"),
--("00000000111111111110000001111111111000"),
--("00000000111111111100000000111111111100"),
--("00000001111111111000000000011111111100"),
--("00000001111111111000000000011111111000"),
--("00000000111111111000000000001111111000"),
--("00000000111111110000000000000111111100"),
--("00000000111111000000000000000011111110"),
--("00000001111110000000000000000001111111"),
--("00000001111111000000000000000001111111"),
--("00000011111111110000000000000001111110"),
--("00000001111111110000000000000000111100")
--);
--constant PinkDead_X_size : integer := 76;
--constant PinkDead_Y_size : integer := 48;
--type PinkDead_color_array is array(0 to PinkDead_Y_size - 1 , 0 to PinkDead_X_size - 1) of std_logic_vector(7 downto 0);
--type PinkDead_bmp_array is array(0 to PinkDead_Y_size - 1 , 0 to PinkDead_X_size - 1) of std_logic;
--constant PinkDead_colors: PinkDead_color_array := (
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F6", x"FA", x"F6", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FA", x"FA", x"F5", x"F5", x"F6", x"F6", x"F5", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F5", x"D1", x"F5", x"FA", x"FA", x"D1", x"D5", x"F5", x"D1", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F6", x"F6", x"F6", x"F5", x"CD", x"AD", x"88", x"60", x"64", x"60", x"60", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B7", x"6D", x"64", x"68", x"68", x"AD", x"D2", x"CE", x"40", x"40", x"40", x"40", x"40", x"40", x"64", x"DF", x"FF", x"FF", x"FB", x"FB", x"FF", x"FF", x"FB", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EA", x"EE", x"EE", x"EE", x"EE", x"E9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"69", x"64", x"40", x"60", x"40", x"40", x"40", x"40", x"D2", x"FB", x"F2", x"EE", x"CE", x"D2", x"F6", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"C9", x"C9", x"C9", x"EE", x"EE", x"E9", x"C9", x"C9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"88", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"69", x"CE", x"60", x"40", x"60", x"40", x"40", x"60", x"C9", x"F2", x"EE", x"F2", x"CE", x"C9", x"C9", x"E9", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"C9", x"C5", x"C9", x"C9", x"C9", x"E9", x"C9", x"C9", x"E9", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FA", x"B1", x"00", x"00", x"00", x"00", x"00", x"49", x"D2", x"F7", x"F6", x"A9", x"40", x"40", x"40", x"40", x"64", x"D2", x"F7", x"F2", x"F2", x"F7", x"CE", x"EE", x"C9", x"C9", x"C9", x"EE", x"E9", x"EE", x"EE", x"C5", x"E9", x"EE", x"EE", x"CD", x"EE", x"C9", x"E9", x"E9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F6", x"D1", x"D1", x"D6", x"DB", x"FA", x"F6", x"D2", x"B2", x"B2", x"AE", x"AE", x"AE", x"F2", x"F7", x"F7", x"F6", x"ED", x"CD", x"D1", x"D1", x"D1", x"D1", x"AD", x"D3", x"F7", x"F7", x"F7", x"F2", x"F7", x"EE", x"EE", x"EE", x"CE", x"C9", x"C9", x"C9", x"C5", x"C9", x"E9", x"E9", x"C9", x"E9", x"C9", x"C9", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"F6", x"D1", x"D2", x"D5", x"D5", x"D1", x"CC", x"F2", x"FB", x"D3", x"F7", x"F7", x"F3", x"F7", x"F7", x"F3", x"F7", x"F7", x"F2", x"CD", x"F5", x"F5", x"F5", x"F1", x"D1", x"89", x"65", x"AD", x"F2", x"F7", x"F2", x"F7", x"F2", x"F2", x"F7", x"F7", x"F2", x"D2", x"F2", x"F2", x"D2", x"F2", x"EE", x"EE", x"EE", x"CE", x"CE", x"EE", x"FB", x"FF", x"FF", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FB", x"D6", x"AD", x"AD", x"AD", x"D1", x"D5", x"D1", x"F6", x"F1", x"F2", x"D2", x"AE", x"AD", x"AD", x"AD", x"D2", x"F6", x"F2", x"F2", x"F2", x"CE", x"F2", x"EE", x"ED", x"CD", x"89", x"20", x"89", x"F7", x"89", x"00", x"69", x"F7", x"F7", x"F7", x"F7", x"F7", x"FB", x"FB", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"D6", x"B1", x"88", x"88", x"6D", x"F5", x"F5", x"D1", x"F1", x"F2", x"D2", x"69", x"8D", x"D5", x"F1", x"F1", x"F6", x"FA", x"FA", x"F6", x"F1", x"CD", x"F2", x"F2", x"F2", x"F2", x"A9", x"00", x"44", x"F7", x"AE", x"00", x"00", x"89", x"C9", x"A9", x"AE", x"AE", x"AE", x"D2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"F1", x"F1", x"D5", x"F6", x"F6", x"F5", x"F1", x"F6", x"F6", x"FB"),
--( x"FF", x"FF", x"FF", x"D6", x"D6", x"A8", x"68", x"88", x"F1", x"AC", x"D1", x"CD", x"CE", x"24", x"48", x"F6", x"FA", x"F6", x"F5", x"FA", x"FA", x"F6", x"F5", x"F1", x"F5", x"F6", x"FA", x"FA", x"F6", x"D1", x"8D", x"8D", x"ED", x"A8", x"40", x"40", x"40", x"60", x"40", x"60", x"40", x"40", x"AD", x"F1", x"F6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"CD", x"CC", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"D1", x"F6"),
--( x"FF", x"FF", x"FF", x"DB", x"D6", x"88", x"84", x"88", x"A8", x"88", x"CD", x"CD", x"CE", x"00", x"68", x"FA", x"FA", x"F5", x"F1", x"F5", x"F6", x"F6", x"F5", x"F6", x"F6", x"F6", x"F6", x"F6", x"FA", x"F6", x"FA", x"FA", x"F5", x"88", x"40", x"60", x"40", x"40", x"60", x"60", x"40", x"40", x"CD", x"F1", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"ED", x"CD", x"F1", x"F5", x"F5", x"F5", x"F1", x"F1", x"D1", x"FB"),
--( x"FF", x"D6", x"AD", x"88", x"AC", x"88", x"84", x"84", x"84", x"84", x"A8", x"EE", x"F2", x"85", x"44", x"B1", x"FA", x"F1", x"CD", x"F5", x"F6", x"F5", x"F5", x"F1", x"F5", x"F5", x"F6", x"F6", x"F6", x"F6", x"F6", x"F5", x"F1", x"84", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"CD", x"CD", x"C9", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"CD", x"D1", x"D6", x"D6", x"D1", x"F1", x"F1", x"F1", x"D1", x"D1", x"FF"),
--( x"FB", x"AC", x"AD", x"AC", x"AC", x"AD", x"88", x"84", x"88", x"88", x"A8", x"CD", x"F2", x"F2", x"AD", x"89", x"89", x"89", x"CD", x"F1", x"F6", x"F6", x"F2", x"F6", x"F6", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F6", x"D2", x"64", x"60", x"60", x"64", x"89", x"A9", x"84", x"AD", x"D1", x"CD", x"D6", x"F7", x"F7", x"F6", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"FB", x"FF", x"FF", x"FB", x"D6", x"F1", x"D1", x"D1", x"FB", x"FF"),
--( x"FF", x"DA", x"FB", x"FF", x"DA", x"DB", x"DA", x"D6", x"DA", x"FB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FB", x"D6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"DB", x"D6", x"D6", x"DA", x"FF", x"FF", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"FB", x"F6", x"F7", x"F6", x"F7", x"FB", x"FF", x"F7", x"F7", x"F7", x"F7", x"FB", x"FF", x"FF", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"FB", x"FF", x"FF")
--);
--constant PinkDead_bmp: PinkDead_bmp_array := (
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000000000000000000000000000000000000000000000000000000"),
--("0000000000000000000000000111111000000000000000000000000000000000000000000000"),
--("0000000000000000000000111111111000000000000000111111111000000000000000000000"),
--("0000000000000000000001111111111100000000000011111111111100000000000000000000"),
--("0000000000000000000111111111111100000000011111111111111110000000000000000000"),
--("0000000000000000011111111111111110011001111111111111111110000000000000000000"),
--("0000000000000000111111111111111111111111111111111111111110000000000000000000"),
--("0000000000000001111111111111111111111111111111111111111100000000000000000000"),
--("0000000001110001111111111111111111111111111111111111111100000000000000000000"),
--("0000000011111111111111111111111111111111111111111111111100000000000000000000"),
--("0000001111111111111111111111111111111111111111111111111100111110000000000000"),
--("0001111111111111111111111111111111111111111111111111111111111111100000000000"),
--("0001111111111111111111111111111111111111111111111111111111111111111111111111"),
--("0001111111111111111111111111111111111111111111111111111111111111111111111111"),
--("0001111111111111111111111111111111111111111111111111111111111111111111111111"),
--("0111111111111111111111111111111111111111111111111111111111111111111111111110"),
--("1111111111111111111111111111111111111111111111111111111111111111111001111110"),
--("0110111111100001110000000111111000111100111000001011111101111100110000001100")
--);
--constant PinkIdle_X_size : integer := 32;
--constant PinkIdle_Y_size : integer := 48;
--type PinkIdle_color_array is array(0 to PinkIdle_Y_size - 1 , 0 to PinkIdle_X_size - 1) of std_logic_vector(7 downto 0);
--type PinkIdle_bmp_array is array(0 to PinkIdle_Y_size - 1 , 0 to PinkIdle_X_size - 1) of std_logic;
--constant PinkIdle_colors: PinkIdle_color_array := (
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"B6", x"B6", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"68", x"64", x"64", x"64", x"64", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"68", x"64", x"64", x"88", x"68", x"88", x"64", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B2", x"64", x"64", x"64", x"88", x"AD", x"D1", x"64", x"68", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"8D", x"64", x"88", x"AD", x"88", x"44", x"44", x"D1", x"AD", x"49", x"B1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"D2", x"D2", x"89", x"A4", x"AD", x"CD", x"B1", x"F6", x"68", x"8D", x"69", x"B6", x"B2", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"D1", x"8D", x"AE", x"D2", x"CE", x"C9", x"C9", x"CD", x"F5", x"CD", x"D1", x"F6", x"D5", x"CD", x"D1", x"DA", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"D6", x"F1", x"F5", x"D5", x"69", x"AE", x"CE", x"CE", x"D2", x"AD", x"F1", x"F6", x"D1", x"AD", x"D1", x"D1", x"AC", x"AD", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"F5", x"F6", x"F6", x"D5", x"69", x"CE", x"C9", x"D2", x"AD", x"AC", x"CD", x"D1", x"D1", x"AD", x"CD", x"AD", x"8D", x"A9", x"CE", x"F2", x"D6", x"D2", x"D2", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"D6", x"D1", x"F5", x"F1", x"D1", x"8D", x"A9", x"CE", x"B2", x"20", x"48", x"88", x"68", x"D1", x"D1", x"CD", x"CE", x"D2", x"CE", x"D2", x"8D", x"49", x"44", x"A9", x"CD", x"FB", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"CD", x"CD", x"F1", x"D1", x"F5", x"F6", x"CD", x"D2", x"65", x"00", x"00", x"40", x"20", x"64", x"D1", x"A8", x"AD", x"CE", x"CE", x"D2", x"85", x"68", x"D5", x"F6", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"F1", x"D1", x"F1", x"D1", x"D1", x"D5", x"D1", x"A9", x"20", x"20", x"40", x"40", x"20", x"20", x"AD", x"D1", x"A9", x"CE", x"D6", x"89", x"48", x"D5", x"F6", x"F5", x"F1", x"AD", x"FB", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"D1", x"F5", x"D5", x"D5", x"D1", x"CD", x"88", x"40", x"40", x"40", x"40", x"20", x"20", x"40", x"D1", x"D1", x"AD", x"D2", x"D7", x"69", x"8D", x"F1", x"D1", x"F1", x"D1", x"AD", x"FB", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"AD", x"CD", x"F6", x"F6", x"D5", x"F5", x"AD", x"20", x"40", x"20", x"20", x"40", x"40", x"44", x"AD", x"AC", x"D1", x"CE", x"D2", x"AE", x"89", x"CD", x"CD", x"CD", x"CD", x"A8", x"D6", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"D6", x"AD", x"D1", x"D5", x"F5", x"F5", x"D1", x"64", x"20", x"20", x"20", x"89", x"CD", x"A9", x"B2", x"D2", x"D6", x"CE", x"CE", x"CE", x"AD", x"CD", x"CD", x"CD", x"D1", x"CD", x"CD", x"FB", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"D1", x"CD", x"F1", x"F1", x"F1", x"CD", x"CD", x"64", x"20", x"89", x"D2", x"CE", x"D2", x"D7", x"D7", x"D2", x"CE", x"CE", x"C9", x"A8", x"D1", x"CD", x"D1", x"F1", x"F1", x"CD", x"D6", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"D6", x"AD", x"CC", x"CD", x"AD", x"A9", x"CD", x"C9", x"64", x"CE", x"CE", x"CE", x"D2", x"D2", x"D2", x"CE", x"CE", x"CE", x"AD", x"AD", x"AD", x"AC", x"A9", x"AD", x"F1", x"D1", x"B1", x"FB", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"D6", x"A9", x"C9", x"C9", x"CE", x"C9", x"C9", x"C9", x"C9", x"CE", x"CE", x"CE", x"CE", x"CE", x"CD", x"AD", x"AD", x"69", x"44", x"20", x"20", x"64", x"CD", x"CC", x"B2", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"CE", x"C9", x"C9", x"CD", x"CD", x"C9", x"C9", x"C9", x"CD", x"CE", x"C9", x"C9", x"CD", x"AD", x"D1", x"D5", x"64", x"20", x"40", x"20", x"64", x"D1", x"AD", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"65", x"64", x"85", x"89", x"89", x"89", x"89", x"85", x"65", x"20", x"69", x"FB", x"B1", x"CD", x"D1", x"88", x"20", x"20", x"20", x"64", x"CD", x"AD", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"85", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"40", x"A9", x"D6", x"B6", x"AD", x"B1", x"D1", x"20", x"20", x"40", x"88", x"AD", x"DB", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"CD", x"64", x"00", x"24", x"20", x"00", x"65", x"85", x"89", x"C9", x"C9", x"C9", x"D2", x"8D", x"AD", x"8D", x"20", x"40", x"88", x"D6", x"DB", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"CE", x"64", x"20", x"CD", x"C9", x"20", x"44", x"EE", x"CE", x"C9", x"C9", x"C9", x"D2", x"DB", x"DB", x"DB", x"DA", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"A9", x"C9", x"A9", x"00", x"44", x"CE", x"C9", x"00", x"20", x"CE", x"CE", x"C9", x"CD", x"A9", x"A9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"AE", x"D2", x"D2", x"A9", x"00", x"44", x"C9", x"C9", x"20", x"00", x"89", x"C9", x"C9", x"CE", x"C9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D2", x"D7", x"D7", x"CE", x"20", x"20", x"A5", x"A9", x"20", x"00", x"89", x"C9", x"CE", x"CE", x"CE", x"CE", x"DF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"F7", x"D2", x"D7", x"D7", x"D7", x"D2", x"24", x"00", x"89", x"CE", x"20", x"20", x"CE", x"CE", x"D2", x"D6", x"D6", x"A9", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FB", x"D2", x"D7", x"D7", x"D7", x"D7", x"D2", x"24", x"40", x"A5", x"CE", x"24", x"64", x"D2", x"D7", x"D7", x"D7", x"D7", x"D2", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"D2", x"D6", x"D7", x"D7", x"D6", x"D7", x"D7", x"AE", x"CE", x"C9", x"A5", x"A9", x"CD", x"D6", x"D7", x"D7", x"D7", x"D7", x"D7", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"CE", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"C9", x"CD", x"D2", x"C9", x"CE", x"D6", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"D2", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"CE", x"C9", x"DB", x"F7", x"C9", x"CE", x"D6", x"D6", x"D7", x"D7", x"D7", x"D7", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"F7", x"D2", x"D7", x"D7", x"D7", x"D3", x"D2", x"D2", x"CE", x"D6", x"FF", x"FB", x"A9", x"CE", x"CE", x"D6", x"D7", x"D7", x"D7", x"D7", x"CE", x"D2", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"D2", x"D2", x"D6", x"D6", x"D7", x"D7", x"D6", x"CE", x"D2", x"FF", x"FF", x"FF", x"D2", x"C9", x"D2", x"D2", x"D2", x"D6", x"D7", x"D7", x"D2", x"D2", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"F2", x"EE", x"EE", x"D2", x"D7", x"D7", x"CE", x"A9", x"FB", x"FF", x"FF", x"FF", x"FF", x"CE", x"D2", x"D7", x"D7", x"D6", x"CE", x"D2", x"D2", x"CE", x"CA", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"CE", x"CE", x"EE", x"EE", x"D2", x"D2", x"CE", x"CD", x"D7", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"D2", x"D7", x"D7", x"D2", x"CE", x"CE", x"CE", x"EE", x"CE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"D7", x"C9", x"EE", x"EE", x"EE", x"CE", x"D2", x"CE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"CE", x"D2", x"CE", x"CE", x"EE", x"CE", x"CE", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"CE", x"CE", x"EE", x"EE", x"EE", x"EE", x"CE", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"CE", x"CE", x"CE", x"EE", x"CE", x"EE", x"CE", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"D2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CD", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"D2", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"D2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"CE", x"EE", x"CE", x"CE", x"EE", x"EE", x"CD", x"D2", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"F7", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"FB", x"FF", x"FF"),
--( x"FF", x"FF", x"F6", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"C9", x"EE", x"EE", x"EE", x"EE", x"F2", x"C9", x"D2", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"F7", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"CD", x"EE", x"EE", x"EE", x"EE", x"CD", x"CD", x"FB", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FB", x"CD", x"CD", x"CD", x"CD", x"D2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D6", x"CE", x"CD", x"CD", x"F1", x"D1", x"D6", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"D6", x"F1", x"F5", x"F1", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F5", x"F5", x"F5", x"D1", x"D6", x"FF"),
--( x"FF", x"FF", x"D6", x"F1", x"F5", x"F1", x"F5", x"F1", x"CC", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F1", x"F1", x"F1", x"F1", x"F1", x"CD", x"DA"),
--( x"D6", x"D1", x"D1", x"D1", x"F1", x"F1", x"F1", x"F1", x"CD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"F5", x"CD", x"D1", x"D1", x"CD", x"CD", x"AD"),
--( x"CC", x"A8", x"CD", x"CD", x"D1", x"D1", x"CD", x"B1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"D2", x"D6", x"D1", x"D1", x"D6", x"DA", x"FB"),
--( x"DA", x"DA", x"DA", x"FB", x"DB", x"FA", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
--);
--constant PinkIdle_bmp: PinkIdle_bmp_array := (
--("00000000000000011111000000000000"),
--("00000000000000111111100000000000"),
--("00000000000000111111110000000000"),
--("00000000000001111111111000000000"),
--("00000000000011111111111100000000"),
--("00000000111111111111111100000000"),
--("00001111111111111111111000000000"),
--("00011111111111111111110000000000"),
--("00111111111111111111111111110000"),
--("00111111111111111111111111110000"),
--("00111111111111111111111111110000"),
--("01111111111111111111111111111000"),
--("01111111111111111111111111111000"),
--("00111111111111111111111111111000"),
--("00111111111111111111111111111100"),
--("00011111111111111111111111111100"),
--("00011111111111111111111111111110"),
--("00001111111111111111111111111110"),
--("00000001111111111111111111111110"),
--("00000000111111111111111111111110"),
--("00000000111111111111111111111110"),
--("00000001111111111111111111111100"),
--("00000001111111111111111111100000"),
--("00000011111111111111111000000000"),
--("00000111111111111111110000000000"),
--("00000111111111111111111000000000"),
--("00001111111111111111111000000000"),
--("00011111111111111111111000000000"),
--("00011111111111111111111000000000"),
--("00111111111111111111111000000000"),
--("00111111111111111111111100000000"),
--("00111111111101111111111110000000"),
--("00111111111000111111111111000000"),
--("00111111111000011111111111000000"),
--("00111111111000011111111111100000"),
--("01111111111000001111111111100000"),
--("01111111111000000111111111110000"),
--("00111111111000000011111111110000"),
--("00111111111000000001111111111000"),
--("00111111111000000001111111111100"),
--("00111111111100000000111111111000"),
--("00111111111000000000011111111100"),
--("00011111110000000000001111111100"),
--("00011111100000000000000011111110"),
--("00111111110000000000000111111111"),
--("11111111110000000000000111111111"),
--("11111111100000000000000111111111"),
--("11111110000000000000000000000000")
--);
--constant PinkWon_X_size : integer := 38;
--constant PinkWon_Y_size : integer := 48;
--type PinkWon_color_array is array(0 to PinkWon_Y_size - 1 , 0 to PinkWon_X_size - 1) of std_logic_vector(7 downto 0);
--type PinkWon_bmp_array is array(0 to PinkWon_Y_size - 1 , 0 to PinkWon_X_size - 1) of std_logic;
--constant PinkWon_colors: PinkWon_color_array := (
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"88", x"88", x"88", x"AC", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"88", x"88", x"88", x"A8", x"88", x"88", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"8D", x"88", x"AD", x"D1", x"AD", x"88", x"84", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"20", x"AD", x"D1", x"89", x"64", x"88", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"AD", x"A8", x"AD", x"CD", x"F1", x"D1", x"D1", x"A8", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"D2", x"D1", x"CD", x"AC", x"AC", x"D5", x"FA", x"F1", x"D1", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"F2", x"CE", x"84", x"88", x"AD", x"CD", x"F1", x"F2", x"F2", x"A9", x"CD", x"FB", x"FB", x"FB", x"FB", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F2", x"D2", x"64", x"20", x"40", x"64", x"64", x"68", x"8D", x"F2", x"F2", x"EE", x"F2", x"F2", x"CE", x"C9", x"CA", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F2", x"F2", x"F3", x"AE", x"00", x"40", x"60", x"40", x"40", x"00", x"8D", x"F2", x"F7", x"F7", x"F7", x"F7", x"89", x"89", x"ED", x"FB", x"FF", x"FF", x"FF", x"DB", x"8D", x"20", x"60", x"D1", x"D5", x"D1", x"D1", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"EE", x"F7", x"8D", x"20", x"40", x"40", x"84", x"64", x"64", x"F2", x"F2", x"F7", x"F7", x"F7", x"AE", x"B1", x"FA", x"F5", x"D1", x"FB", x"FF", x"FF", x"69", x"64", x"88", x"84", x"A8", x"AD", x"D1", x"D6", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"A8", x"EE", x"F7", x"AE", x"40", x"40", x"40", x"20", x"40", x"D2", x"F7", x"D2", x"F2", x"F2", x"CE", x"A9", x"F6", x"FA", x"F6", x"F1", x"F6", x"FF", x"8D", x"40", x"D1", x"F5", x"C8", x"A8", x"DB", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CC", x"EE", x"F3", x"CD", x"60", x"40", x"40", x"00", x"8D", x"F7", x"F7", x"F2", x"F2", x"EE", x"A9", x"D1", x"FA", x"FA", x"F6", x"F5", x"F1", x"AD", x"40", x"60", x"64", x"64", x"D1", x"DA", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"CD", x"CD", x"F1", x"D1", x"A9", x"40", x"44", x"F7", x"F7", x"F3", x"F7", x"F2", x"EE", x"C9", x"F1", x"F5", x"F6", x"FA", x"F5", x"CC", x"20", x"20", x"40", x"00", x"8D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CC", x"A8", x"CD", x"F5", x"F6", x"F1", x"84", x"AE", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"C9", x"CD", x"F1", x"F1", x"F1", x"D1", x"CD", x"A8", x"60", x"20", x"44", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"CC", x"C8", x"F1", x"F6", x"F5", x"CC", x"AD", x"F7", x"F7", x"F7", x"F6", x"EE", x"EE", x"EE", x"CD", x"AD", x"F1", x"F1", x"CD", x"CD", x"F1", x"F5", x"D1", x"84", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"A8", x"CC", x"F1", x"F1", x"CD", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"CD", x"CD", x"CD", x"F5", x"F5", x"F5", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D6", x"AD", x"A8", x"CD", x"F2", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"D2", x"D6", x"D1", x"F5", x"F5", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"FF", x"FF", x"D6", x"CD", x"CD", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"60", x"85", x"CD", x"EE", x"EE", x"EE", x"EE", x"A9", x"65", x"40", x"64", x"DB", x"FF", x"FF", x"FF", x"D6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"44", x"00", x"20", x"40", x"20", x"20", x"20", x"00", x"20", x"65", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"CE", x"00", x"20", x"65", x"00", x"00", x"65", x"A9", x"CE", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"89", x"00", x"89", x"EE", x"64", x"20", x"CE", x"F2", x"F2", x"EE", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EA", x"24", x"00", x"CE", x"EE", x"A9", x"00", x"A9", x"F2", x"EE", x"EA", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"20", x"20", x"EE", x"F2", x"C9", x"00", x"69", x"EE", x"EE", x"F2", x"F2", x"F2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"D2", x"20", x"44", x"EE", x"EE", x"CE", x"00", x"65", x"EE", x"F7", x"F7", x"F7", x"F7", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F7", x"8D", x"00", x"44", x"F2", x"EE", x"CE", x"00", x"65", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"F7", x"69", x"20", x"AE", x"F2", x"EE", x"C9", x"20", x"69", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"D7", x"B2", x"D2", x"F7", x"F2", x"EE", x"C9", x"64", x"A9", x"F2", x"F7", x"F7", x"D7", x"F7", x"F2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"F7", x"F7", x"FB", x"F7", x"F2", x"EE", x"E9", x"C9", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"F7", x"D7", x"D7", x"F3", x"F2", x"EE", x"C9", x"D6", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"CE", x"FF", x"F6", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F7", x"FB", x"F7", x"F2", x"EE", x"E9", x"F2", x"FF", x"FB", x"EE", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"FB", x"FF", x"FF", x"F2", x"F2", x"F2", x"D7", x"F7", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C5", x"EE", x"EE", x"EE", x"EE", x"E9", x"C9", x"FB", x"FF", x"FF", x"F6", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"E9", x"E9", x"E9", x"EE", x"EE", x"E9", x"C9", x"FB", x"FF", x"FF", x"FF", x"CE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"EE", x"EE", x"CE", x"EE", x"EE", x"E9", x"CE", x"FB", x"FF", x"FF", x"FF", x"D2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"D2", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"E9", x"EE", x"EE", x"ED", x"EE", x"EE", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"E9", x"EE", x"EE", x"EE", x"EE", x"E9", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"D2", x"C5", x"E9", x"EE", x"CA", x"EA", x"EE", x"C9", x"C5", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FB", x"D2", x"E9", x"C9", x"C9", x"E9", x"C9", x"C9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"EE", x"ED", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"ED", x"CD", x"CD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"D6", x"CD", x"ED", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"F1", x"CC", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F5", x"F1", x"D1", x"CD", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F1", x"F1", x"ED", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"F1", x"F5", x"F5", x"F1", x"CC", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"CD", x"F1", x"F5", x"F1", x"F5", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"D6", x"D1", x"F1", x"F1", x"F5", x"F1", x"CC", x"C8", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"ED", x"F1", x"F1", x"F1", x"F1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"D6", x"CD", x"CD", x"D1", x"D1", x"F1", x"F1", x"D1", x"B1", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"F1", x"F1", x"D1", x"F1", x"CD", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"D6", x"DA", x"FA", x"FA", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"D1", x"D1", x"D1", x"A8", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
--);
--constant PinkWon_bmp: PinkWon_bmp_array := (
--("00000000000111111000000000000000000000"),
--("00000000001111111100000000000000000000"),
--("00000000001111111100000000000000000000"),
--("00000000001111111100000000000000000000"),
--("00000000011111111110000000000000000000"),
--("00000001111111111111000000000000000000"),
--("00000001111111111111111111000000000000"),
--("00000011111111111111111111000001100000"),
--("00000111111111111111111111000111111110"),
--("00000111111111111111111111100111111110"),
--("00000111111111111111111111101111111000"),
--("00000111111111111111111111111111110000"),
--("00000111111111111111111111111111100000"),
--("00000111111111111111111111111110000000"),
--("00000111111111111111111111111110000000"),
--("00000011111111111111111111111100000000"),
--("00000011111111111111111111111000000000"),
--("00000000111111111111110011111000000000"),
--("00000000011111111111110001100000000000"),
--("00000000011111111111100000000000000000"),
--("00000000111111111111110000000000000000"),
--("00000000111111111111110000000000000000"),
--("00000000111111111111111000000000000000"),
--("00000000111111111111111000000000000000"),
--("00000001111111111111111000000000000000"),
--("00000001111111111111111000000000000000"),
--("00000011111111111111111100000000000000"),
--("00000011111111111111111100000000000000"),
--("00000011111111111111111100000000000000"),
--("00000011111111111111111100000000000000"),
--("00000011111111101111111100000000000000"),
--("00000011111111101111111110000000000000"),
--("00000011111111100111111110000000000000"),
--("00000011111111100111111111000000000000"),
--("00000111111111100011111111000000000000"),
--("00000111111111100011111111100000000000"),
--("00000111111111000011111111100000000000"),
--("00000111111111000001111111100000000000"),
--("00001111111111000001111111110000000000"),
--("00001111111111000001111111110000000000"),
--("00001111111110000000111111100000000000"),
--("00000011111100000000111111000000000000"),
--("00000011111000000000001111100000000000"),
--("00000111111100000000001111110000000000"),
--("00001111111100000000001111110000000000"),
--("00111111111100000000001111111000000000"),
--("01111111111100000000001111111110000000"),
--("01111111000000000000000111111110000000")
--);
--constant PinkPunch_X_size : integer := 44;
--constant PinkPunch_Y_size : integer := 48;
--type PinkPunch_color_array is array(0 to PinkPunch_Y_size - 1 , 0 to PinkPunch_X_size - 1) of std_logic_vector(7 downto 0);
--type PinkPunch_bmp_array is array(0 to PinkPunch_Y_size - 1 , 0 to PinkPunch_X_size - 1) of std_logic;
--constant PinkPunch_colors: PinkPunch_color_array := (
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"B2", x"8D", x"B2", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"88", x"88", x"88", x"88", x"B1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"68", x"40", x"40", x"40", x"69", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"84", x"88", x"88", x"88", x"88", x"68", x"AC", x"FB", x"FF", x"FF", x"FF", x"FF", x"F6", x"64", x"40", x"60", x"60", x"40", x"B2", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"8C", x"84", x"88", x"AC", x"AD", x"D1", x"AC", x"84", x"D6", x"FF", x"FF", x"FF", x"FF", x"D1", x"D1", x"8D", x"40", x"40", x"40", x"65", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"88", x"AC", x"A8", x"88", x"24", x"8D", x"F6", x"CD", x"D6", x"DA", x"FF", x"FF", x"FF", x"D6", x"F5", x"88", x"40", x"60", x"40", x"40", x"DB"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"AD", x"AC", x"88", x"88", x"A4", x"D1", x"F1", x"D5", x"AD", x"44", x"88", x"F6", x"FB", x"D6", x"FF", x"FF", x"FF", x"FF", x"FA", x"64", x"40", x"60", x"40", x"40", x"D6"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"B2", x"88", x"88", x"88", x"88", x"88", x"D1", x"F5", x"F1", x"F6", x"FA", x"F1", x"D1", x"FA", x"FB", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"69", x"AD", x"F6", x"CD", x"60", x"D7"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"EE", x"88", x"88", x"88", x"88", x"D1", x"F1", x"F5", x"FA", x"FA", x"F1", x"CD", x"AD", x"D6", x"F6", x"F6", x"F6", x"FB", x"FF", x"FB", x"FF", x"FF", x"FF", x"D1", x"F6", x"FA", x"F6", x"CD", x"DA"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"EE", x"CD", x"64", x"88", x"CC", x"D1", x"F6", x"FA", x"FA", x"FA", x"F6", x"F5", x"F1", x"F1", x"F5", x"F6", x"F6", x"F6", x"F1", x"D1", x"D1", x"D1", x"D6", x"D6", x"FA", x"F6", x"F5", x"FA", x"F1", x"FA"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"EE", x"F2", x"CE", x"88", x"A9", x"F1", x"F1", x"F6", x"FA", x"F6", x"F5", x"F5", x"F5", x"F6", x"FA", x"FA", x"FA", x"F6", x"F6", x"F6", x"F5", x"F1", x"F6", x"F5", x"F6", x"FA", x"F5", x"F1", x"FA", x"F5", x"F6"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"EE", x"EE", x"F2", x"A9", x"D2", x"F2", x"F1", x"FA", x"F6", x"F5", x"F6", x"FA", x"F6", x"F6", x"F6", x"FA", x"F6", x"F6", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"FA"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"EE", x"F2", x"F7", x"D2", x"D6", x"F2", x"F1", x"FA", x"F6", x"F5", x"F6", x"FA", x"FA", x"F5", x"F1", x"F1", x"F1", x"F6", x"F5", x"F6", x"F6", x"F5", x"F5", x"F6", x"F5", x"F5", x"F5", x"F5", x"D1", x"D1", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F1", x"EE", x"EE", x"EE", x"F7", x"F2", x"F2", x"D7", x"F6", x"F6", x"FA", x"F5", x"F6", x"F6", x"F5", x"F1", x"F1", x"AC", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"CD", x"F1", x"F1", x"D1", x"F5", x"F1", x"B1", x"FB", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F1", x"E9", x"EE", x"F6", x"F7", x"F2", x"F7", x"F7", x"D2", x"D1", x"D5", x"FA", x"FA", x"F6", x"F5", x"F1", x"A8", x"AC", x"AD", x"CD", x"CD", x"D1", x"D1", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"ED", x"F5", x"F1", x"C9", x"EE", x"F2", x"F2", x"F2", x"EE", x"F7", x"D2", x"69", x"24", x"68", x"8D", x"D1", x"CD", x"68", x"44", x"69", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"F5", x"ED", x"E9", x"F2", x"F2", x"EE", x"EE", x"F2", x"F3", x"F7", x"B2", x"45", x"00", x"20", x"00", x"00", x"00", x"00", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"F1", x"F1", x"C9", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F3", x"F2", x"D6", x"B2", x"24", x"00", x"00", x"00", x"00", x"48", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"AD", x"CD", x"C9", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"A9", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"C9", x"C9", x"C9", x"A9", x"C9", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"89", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"89", x"85", x"89", x"89", x"A5", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"89", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"EE", x"F2", x"F7", x"F7", x"CE", x"C9", x"C9", x"EE", x"EE", x"EE", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F6", x"F2", x"F2", x"EE", x"C9", x"C9", x"C5", x"C5", x"C5", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F7", x"F7", x"F2", x"EE", x"EE", x"40", x"44", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"F2", x"D2", x"F7", x"F7", x"F7", x"F7", x"EE", x"CE", x"24", x"44", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"EE", x"EE", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"C9", x"20", x"45", x"F3", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"C9", x"EE", x"F6", x"F7", x"F7", x"D7", x"F7", x"F7", x"EE", x"84", x"00", x"45", x"F2", x"F2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"E9", x"84", x"00", x"85", x"F2", x"F2", x"F2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"EE", x"C5", x"85", x"00", x"C9", x"F2", x"F2", x"F2", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"E9", x"C5", x"C9", x"C9", x"CE", x"EE", x"EE", x"EE", x"F2", x"F6", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F2", x"F6", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"CE", x"C5", x"C9", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F6", x"F6", x"C9", x"C5", x"C9", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"D2", x"F2", x"FF", x"FF", x"FB", x"CE", x"C9", x"E9", x"C9", x"E9", x"EE", x"EE", x"EE", x"EE", x"E9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C5", x"E9", x"C9", x"E9", x"CE", x"EE", x"EE", x"E9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"F3", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"EE", x"EA", x"EE", x"EE", x"EE", x"EE", x"E9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"E9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"E9", x"EE", x"EE", x"CD", x"E9", x"EE", x"EE", x"E9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F7", x"F7", x"F6", x"F2", x"F2", x"F2", x"EE", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"EE", x"EA", x"EE", x"EE", x"E9", x"E9", x"E9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"F6", x"E9", x"F2", x"F6", x"F3", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"C9", x"EE", x"CE", x"ED", x"EE", x"C9", x"E9", x"E9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"D2", x"A4", x"CD", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"EE", x"EE", x"EE", x"E9", x"C9", x"EE", x"E9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"D2", x"CC", x"CD", x"CD", x"EE", x"F2", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"EE", x"E9", x"EE", x"C9", x"C9", x"EE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"D6", x"D1", x"F5", x"F1", x"F1", x"D1", x"CD", x"C9", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"EE", x"EE", x"C9", x"C9", x"C9", x"C9", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FB", x"D1", x"F1", x"F1", x"F5", x"F1", x"D1", x"D2", x"D2", x"E9", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"CD", x"C9", x"CD", x"F7", x"F2", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"D1", x"F1", x"F5", x"F5", x"F1", x"CD", x"FB", x"FF", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"CC", x"F1", x"CD", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"F1", x"F1", x"F5", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"CD", x"D1", x"F1", x"D1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"F6", x"F1", x"F5", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"ED", x"F1", x"F1", x"F1", x"ED", x"F1", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"F1", x"F1", x"F5", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"CC", x"CC", x"CD", x"ED", x"CC", x"ED", x"ED", x"D1", x"CD", x"D1", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FA", x"CD", x"F5", x"F5", x"F1", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D2", x"D2", x"B1", x"D2", x"D6", x"D1", x"CD", x"CD", x"D1", x"CD", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"D6", x"F1", x"D1", x"CD", x"D1", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
--);
--constant PinkPunch_bmp: PinkPunch_bmp_array := (
--("00000000000000000000000000000000000000000000"),
--("00000000000000000000000001111000000001111000"),
--("00000000000000000000000011111110000011111100"),
--("00000000000000000000000111111111000011111110"),
--("00000000000000000000000111111111000011111110"),
--("00000000000000000000001111111111100011111111"),
--("00000000000000000011111111111111100001111111"),
--("00000000000000001111111111111111100000111111"),
--("00000000000001111111111111111111101000111111"),
--("00000000000011111111111111111111111111111111"),
--("00000000000111111111111111111111111111111111"),
--("00000000000111111111111111111111111111111111"),
--("00000000000111111111111111111111111111111110"),
--("00000000001111111111111111111111111111111110"),
--("00000000001111111111111111111111111110000000"),
--("00000000011111111111111111111110000000000000"),
--("00000000011111111111111111111111000000000000"),
--("00000000011111111111111111111111100000000000"),
--("00000000001111111111111111111111000000000000"),
--("00000000000000111111111111111111000000000000"),
--("00000000000000011111111111111110000000000000"),
--("00000000000000111111111111111000000000000000"),
--("00000000000001111111111111111000000000000000"),
--("00000000000001111111111111110000000000000000"),
--("00000000000011111111111111111000000000000000"),
--("00000000000001111111111111111100000000000000"),
--("00000000000001111111111111111100000000000000"),
--("00000000000001111111111111111110000000000000"),
--("00000000000011111111111111111111000000000000"),
--("00000000000111111111111111111111100000000000"),
--("00000000000111111111111111111111110000000000"),
--("00000000001111111111111111111111111000000000"),
--("00000000011111111111100111111111111000000000"),
--("00000000111111111111000001111111111000000000"),
--("00000001111111111110000001111111111000000000"),
--("00000011111111111100000001111111111000000000"),
--("00000111111111111000000001111111111000000000"),
--("00001111111111110000000001111111111000000000"),
--("00001111111111100000000001111111111000000000"),
--("00001111111111000000000001111111111000000000"),
--("01111111111110000000000001111111111000000000"),
--("11111111111100000000000000111111111000000000"),
--("01111111011000000000000000111110000000000000"),
--("00111110000000000000000001111111000000000000"),
--("00111110000000000000000001111111110000000000"),
--("00111100000000000000000011111111111110000000"),
--("01111111000000000000000001111111111111000000"),
--("00111111000000000000000000000000000000000000")
--);
--constant PinkShoot_X_size : integer := 54;
--constant PinkShoot_Y_size : integer := 48;
--type PinkShoot_color_array is array(0 to PinkShoot_Y_size - 1 , 0 to PinkShoot_X_size - 1) of std_logic_vector(7 downto 0);
--type PinkShoot_bmp_array is array(0 to PinkShoot_Y_size - 1 , 0 to PinkShoot_X_size - 1) of std_logic;
--constant PinkShoot_colors: PinkShoot_color_array := (
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D6", x"D6", x"D2", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"88", x"88", x"84", x"84", x"88", x"AC", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"A8", x"84", x"88", x"A8", x"AC", x"AC", x"88", x"88", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F5", x"FB", x"FA", x"F6", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"88", x"88", x"88", x"D1", x"6D", x"8D", x"D1", x"AC", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D1", x"B1", x"F5", x"D6", x"F6", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B1", x"B1", x"AD", x"A8", x"D1", x"AC", x"F1", x"8D", x"24", x"D5", x"F6", x"D6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"AD", x"60", x"40", x"64", x"AD", x"F1", x"FA", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AD", x"88", x"88", x"84", x"84", x"CD", x"D1", x"F5", x"F6", x"F6", x"AD", x"D1", x"FF", x"D6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"A8", x"40", x"40", x"40", x"40", x"60", x"CD", x"F6", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F6", x"8C", x"88", x"88", x"88", x"AD", x"CD", x"CE", x"F6", x"D7", x"F2", x"F6", x"F2", x"F6", x"D6", x"AE", x"A9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FA", x"F6", x"FA", x"FA", x"FA", x"AD", x"88", x"60", x"40", x"40", x"20", x"8D", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"EE", x"A9", x"64", x"88", x"AD", x"D2", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F3", x"AE", x"44", x"AD", x"CD", x"CD", x"F2", x"F6", x"F6", x"D6", x"FB", x"F6", x"F6", x"F5", x"F6", x"F6", x"F5", x"F6", x"FA", x"FA", x"84", x"40", x"20", x"89", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"EE", x"F2", x"AD", x"88", x"CE", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F7", x"F2", x"AD", x"24", x"D1", x"FA", x"F6", x"F5", x"F1", x"F1", x"F5", x"F5", x"F5", x"FA", x"F6", x"F6", x"FA", x"FA", x"F6", x"F6", x"F5", x"D1", x"60", x"40", x"B2", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"EE", x"CD", x"AD", x"CE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F3", x"F7", x"F2", x"A9", x"20", x"68", x"F5", x"F5", x"F6", x"FA", x"F6", x"F6", x"F6", x"F6", x"F6", x"F1", x"F5", x"F6", x"F5", x"F6", x"F5", x"ED", x"CD", x"D2", x"B2", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"F2", x"F2", x"AD", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"AD", x"20", x"AD", x"F5", x"F6", x"FA", x"FA", x"FA", x"F6", x"F6", x"F6", x"F6", x"F6", x"F5", x"F5", x"F1", x"CD", x"CD", x"D6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"EE", x"EE", x"F2", x"F7", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D2", x"20", x"24", x"ED", x"F1", x"F5", x"F1", x"F1", x"F1", x"F1", x"F1", x"D1", x"D1", x"D1", x"D1", x"AD", x"AD", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"EE", x"EA", x"EE", x"F7", x"F3", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"69", x"24", x"CD", x"ED", x"F1", x"D1", x"CD", x"CD", x"CD", x"D1", x"D6", x"D6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F5", x"F1", x"C9", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"D7", x"F2", x"F7", x"65", x"00", x"AC", x"AC", x"64", x"A4", x"AD", x"DA", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F5", x"F5", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"CE", x"65", x"20", x"64", x"A5", x"CE", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F1", x"F5", x"ED", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"C9", x"E9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D1", x"CD", x"CC", x"C8", x"C9", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"CE", x"CE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D6", x"D6", x"D6", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"85", x"85", x"85", x"85", x"85", x"A9", x"CD", x"C9", x"89", x"65", x"65", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"CE", x"C9", x"CE", x"CE", x"D2", x"CE", x"A9", x"69", x"24", x"20", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F7", x"F7", x"F2", x"F2", x"EE", x"F2", x"A9", x"44", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"F2", x"EE", x"EE", x"CE", x"20", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"F2", x"EE", x"F2", x"F2", x"D2", x"F7", x"F7", x"F7", x"F6", x"EE", x"AD", x"00", x"89", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F2", x"D7", x"F7", x"F7", x"F7", x"F7", x"EE", x"A9", x"00", x"89", x"F2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C5", x"C9", x"CE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"EE", x"64", x"00", x"AD", x"F7", x"D6", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"C9", x"40", x"00", x"A9", x"F2", x"F2", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"EE", x"C5", x"20", x"20", x"EE", x"F2", x"F2", x"F3", x"D7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"C9", x"C5", x"A5", x"85", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"C5", x"C9", x"E9", x"EA", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"F2", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"D2", x"CE", x"C5", x"C5", x"C9", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"D6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D2", x"F2", x"FF", x"FB", x"CD", x"C5", x"E9", x"E9", x"EE", x"E9", x"E9", x"EE", x"EE", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"C9", x"C9", x"E9", x"ED", x"EE", x"ED", x"EE", x"EA", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"C9", x"EA", x"EE", x"EE", x"CD", x"EE", x"ED", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"E9", x"E9", x"EE", x"CD", x"EE", x"EE", x"EE", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"EE", x"F2", x"D7", x"F7", x"F2", x"F2", x"EE", x"EE", x"E9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"E9", x"EE", x"EE", x"ED", x"EE", x"C9", x"EA", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"F2", x"F7", x"F7", x"F3", x"F2", x"F2", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"E9", x"EE", x"EE", x"EE", x"EE", x"C9", x"E9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"ED", x"A5", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"E9", x"EE", x"EE", x"CE", x"E9", x"E9", x"E9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FF", x"FF", x"CD", x"A8", x"CD", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"EE", x"EE", x"EE", x"C9", x"C9", x"E9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"F6", x"F6", x"F1", x"F1", x"CD", x"CD", x"EE", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"E9", x"EE", x"EE", x"C9", x"C5", x"C9", x"E9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FB", x"D1", x"F1", x"F1", x"F1", x"F1", x"F1", x"CD", x"C9", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"E9", x"C9", x"C9", x"C9", x"CE", x"C9", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FA", x"F1", x"F5", x"F5", x"F5", x"F1", x"CD", x"FB", x"FB", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"D1", x"AC", x"D6", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"D2", x"F1", x"F5", x"F5", x"F1", x"D6", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"F1", x"D1", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"CD", x"F5", x"F5", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"CD", x"CD", x"F1", x"F1", x"F1", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"D1", x"F5", x"F5", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"EC", x"F1", x"ED", x"F1", x"ED", x"F1", x"F1", x"ED", x"D1", x"D6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"F1", x"F5", x"F5", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"AD", x"AD", x"AC", x"CD", x"D1", x"D1", x"CD", x"CD", x"CD", x"F1", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FB", x"F1", x"F1", x"D1", x"D1", x"D5", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"FF", x"FB", x"FA", x"DA", x"DB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
--( x"FF", x"FF", x"FB", x"F6", x"DA", x"D6", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
--);
--constant PinkShoot_bmp: PinkShoot_bmp_array := (
--("000000000000000000000000000000000000000000000000000000"),
--("000000000000000000000000111110000000000000000000000000"),
--("000000000000000000000001111111100000000000000000000000"),
--("000000000000000000000001111111110000000000000001111000"),
--("000000000000000000000011111111110000000000000011111100"),
--("000000000000000000011111111111111000000000000111111110"),
--("000000000000000001111111111111011000000000001111111110"),
--("000000000000001111111111111111111000000111111111111100"),
--("000000000000111111111111111111111111111111111111111000"),
--("000000000001111111111111111111111111111111111111110000"),
--("000000000001111111111111111111111111111111111111100000"),
--("000000000001111111111111111111111111111111111100000000"),
--("000000000011111111111111111111111111111111110000000000"),
--("000000000011111111111111111111111111111000000000000000"),
--("000000000111111111111111111111111110000000000000000000"),
--("000000000111111111111111111111111000000000000000000000"),
--("000000000111111111111111111111110000000000000000000000"),
--("000000000111111111111111111111100000000000000000000000"),
--("000000000011111111111111111100000000000000000000000000"),
--("000000000000000111111111111100000000000000000000000000"),
--("000000000000001111111111111000000000000000000000000000"),
--("000000000000011111111111111000000000000000000000000000"),
--("000000000000011111111111111100000000000000000000000000"),
--("000000000000111111111111111100000000000000000000000000"),
--("000000000000111111111111111110000000000000000000000000"),
--("000000000000011111111111111111000000000000000000000000"),
--("000000000000011111111111111111100000000000000000000000"),
--("000000000000111111111111111111110000000000000000000000"),
--("000000000001111111111111111111111000000000000000000000"),
--("000000000001111111111111111111111100000000000000000000"),
--("000000000011111111111111111111111100000000000000000000"),
--("000000000111111111111011111111111110000000000000000000"),
--("000000001111111111110000111111111110000000000000000000"),
--("000000011111111111110000111111111110000000000000000000"),
--("000000111111111111100000111111111110000000000000000000"),
--("000001111111111110000000011111111110000000000000000000"),
--("000011111111111100000000011111111100000000000000000000"),
--("000011111111111000000000011111111100000000000000000000"),
--("000011111111110000000000011111111100000000000000000000"),
--("011111111111100000000000011111111100000000000000000000"),
--("111111111111000000000000011111111100000000000000000000"),
--("111111111110000000000000001111101000000000000000000000"),
--("011111100100000000000000001111110000000000000000000000"),
--("011111100000000000000000111111111000000000000000000000"),
--("011111000000000000000000111111111111000000000000000000"),
--("011111100000000000000000111111111111100000000000000000"),
--("011111110000000000000000001110111111000000000000000000"),
--("001111110000000000000000000000000000000000000000000000")
--);
--
--end player_renderer_package;