library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;
use ieee.std_logic_arith.all;

library lab_project;
use lab_project.STREET_FIGHTER_PCKG.all;

entity player_renderer is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		PlayerState		: in std_logic_vector(2 downto 0);
		player_direction : in std_logic;
		
		is_game_over : in std_logic;
		player_won : in std_logic;
		
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end player_renderer;

architecture behav of player_renderer is 

--constant object_X_size : integer := 26;
--constant object_Y_size : integer := 26;
--constant R_high		: integer := 7;
--constant R_low		: integer := 5;
--constant G_high		: integer := 4;
--constant G_low		: integer := 2;
--constant B_high		: integer := 1;
--constant B_low		: integer := 0;

--type ram_array is array(0 to player_length_t - 1 , 0 to player_width_t - 1) of std_logic_vector(7 downto 0);
--type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;

constant PinkKick_X_size : integer := 84;
constant PinkKick_Y_size : integer := 83;
type PinkKick_color_array is array(0 to PinkKick_Y_size - 1 , 0 to PinkKick_X_size - 1) of std_logic_vector(7 downto 0);
type PinkKick_bmp_array is array(0 to PinkKick_Y_size - 1 , 0 to PinkKick_X_size - 1) of std_logic;
constant PinkKick_colors: PinkKick_color_array := (
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"DA", x"DA", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"D6", x"B1", x"B1", x"B1", x"B1", x"D6", x"D6", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"AD", x"84", x"84", x"84", x"8C", x"D6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FB", x"B1", x"D2", x"D6", x"FB", x"B1", x"B1", x"D1", x"88", x"84", x"88", x"B1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"B1", x"88", x"88", x"88", x"88", x"84", x"84", x"84", x"88", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"B1", x"8C", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"FF", x"FF", x"FF", x"FF", x"D6", x"88", x"88", x"84", x"84", x"88", x"88", x"88", x"A8", x"88", x"84", x"88", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"B6", x"88", x"88", x"88", x"88", x"A8", x"CC", x"AC", x"AC", x"88", x"88", x"88", x"AC", x"CD", x"88", x"88", x"88", x"84", x"84", x"88", x"88", x"88", x"88", x"84", x"88", x"A8", x"88", x"84", x"AC", x"FF", x"FF", x"FF", x"89", x"44", x"88", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"D6", x"88", x"88", x"A8", x"A8", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"A4", x"A8", x"88", x"88", x"88", x"88", x"88", x"88", x"A8", x"A8", x"A8", x"EE", x"A9", x"A8", x"C9", x"C9", x"AD", x"FB", x"8D", x"40", x"64", x"A8", x"F5", x"AD", x"D6", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"88", x"88", x"88", x"88", x"B1", x"B1", x"AC", x"84", x"88", x"D2", x"D6", x"D6", x"D6", x"D6", x"C9", x"64", x"84", x"64", x"84", x"84", x"64", x"A8", x"CE", x"EE", x"85", x"AD", x"F2", x"ED", x"F2", x"C9", x"88", x"84", x"A8", x"AC", x"CD", x"AC", x"F6", x"A8", x"A8", x"AC", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"B1", x"88", x"AC", x"D6", x"FB", x"FF", x"FB", x"AD", x"B1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"D1", x"D1", x"D1", x"D1", x"CC", x"C9", x"D2", x"F2", x"89", x"8D", x"B1", x"F6", x"F5", x"F6", x"F5", x"CD", x"A8", x"ED", x"F5", x"A8", x"A8", x"AD", x"AC", x"AC", x"FA", x"CD", x"A8", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"88", x"AC", x"D6", x"FF", x"FF", x"FF", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F6", x"F7", x"F6", x"F2", x"F2", x"EE", x"F2", x"89", x"44", x"AD", x"F6", x"FA", x"FA", x"FA", x"FA", x"FA", x"F5", x"F1", x"CD", x"AC", x"AC", x"CD", x"AC", x"AD", x"CD", x"F1", x"A8", x"D1", x"A8", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"88", x"D6", x"FF", x"FF", x"FF", x"DA", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"F7", x"FB", x"F7", x"F2", x"F2", x"F2", x"F3", x"F2", x"EE", x"89", x"00", x"8D", x"F6", x"FA", x"FA", x"F6", x"F6", x"FA", x"FA", x"FA", x"F5", x"CD", x"AD", x"44", x"AD", x"CD", x"CD", x"CD", x"AD", x"CD", x"CC", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"AD", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"AD", x"D6", x"FF", x"FF", x"FF", x"D6", x"FF", x"FF", x"FB", x"FB", x"F2", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"AE", x"20", x"00", x"B1", x"FA", x"F1", x"F5", x"F5", x"F5", x"F6", x"F6", x"F6", x"F5", x"D1", x"CD", x"AD", x"24", x"44", x"A8", x"B1", x"FB", x"D1", x"F6", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F5", x"CD", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"D6", x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"F7", x"EE", x"C9", x"EE", x"D2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"CD", x"00", x"00", x"B1", x"F1", x"F1", x"F5", x"F6", x"F5", x"F5", x"F5", x"F1", x"F1", x"F6", x"F1", x"CD", x"AD", x"24", x"6E", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"F1", x"F1", x"CD", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"B2", x"00", x"00", x"8D", x"F1", x"F5", x"F6", x"FA", x"FA", x"FA", x"F6", x"F5", x"F6", x"F6", x"F6", x"CD", x"CD", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"F5", x"F1", x"D1", x"FA", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F7", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"CE", x"64", x"00", x"A8", x"CD", x"F1", x"F6", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F5", x"F1", x"F1", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"F5", x"F5", x"F5", x"D6", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F7", x"F7", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"EE", x"F2", x"A5", x"00", x"88", x"AD", x"F1", x"F5", x"F5", x"F6", x"FA", x"FA", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F5", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F5", x"F5", x"F5", x"F1", x"D2", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F7", x"D2", x"64", x"00", x"68", x"D1", x"F1", x"F5", x"F6", x"F6", x"F5", x"F5", x"F6", x"FA", x"FA", x"FA", x"F6", x"FA", x"F6", x"F5", x"F1", x"D1", x"D6", x"68", x"40", x"40", x"40", x"40", x"B1", x"64", x"60", x"60", x"60", x"40", x"40", x"D1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F5", x"F5", x"F1", x"F1", x"F1", x"D6", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F2", x"F7", x"F7", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"F2", x"A9", x"20", x"00", x"68", x"CD", x"F1", x"F5", x"F1", x"F6", x"F1", x"F1", x"F1", x"F6", x"F6", x"F6", x"FA", x"FA", x"FA", x"FA", x"F1", x"84", x"60", x"60", x"60", x"60", x"60", x"40", x"40", x"40", x"60", x"60", x"60", x"40", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"AC", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"D7", x"F7", x"F2", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F2", x"EE", x"A5", x"00", x"00", x"44", x"88", x"D1", x"F1", x"F6", x"F6", x"F5", x"F1", x"F5", x"F6", x"FA", x"FA", x"FA", x"F6", x"F6", x"AD", x"40", x"60", x"60", x"40", x"60", x"40", x"40", x"60", x"40", x"60", x"60", x"60", x"40", x"D1", x"D1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"A8", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"F7", x"F7", x"F7", x"EE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F2", x"F2", x"F3", x"A9", x"89", x"00", x"20", x"89", x"D1", x"F5", x"FA", x"FA", x"F6", x"F6", x"FA", x"FA", x"FA", x"F6", x"F6", x"F6", x"AD", x"40", x"40", x"60", x"60", x"40", x"40", x"40", x"60", x"60", x"60", x"60", x"40", x"40", x"D1", x"F1", x"CC", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"F5", x"F1", x"F5", x"F5", x"F5", x"F1", x"CC", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"F7", x"D7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F7", x"F7", x"F2", x"F7", x"F3", x"CE", x"CD", x"C9", x"C9", x"AD", x"D1", x"F1", x"F1", x"F1", x"F1", x"F5", x"F5", x"F1", x"F1", x"F1", x"A8", x"60", x"60", x"60", x"60", x"40", x"40", x"40", x"60", x"60", x"60", x"40", x"40", x"40", x"D1", x"CD", x"CD", x"DB", x"FF", x"FB", x"FB", x"F7", x"F7", x"F7", x"F7", x"FB", x"D6", x"CD", x"F1", x"F1", x"F5", x"F1", x"F1", x"F5", x"F5", x"F5", x"F1", x"DA", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"F2", x"F7", x"F7", x"F7", x"EE", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"EE", x"F2", x"F7", x"F7", x"F2", x"EE", x"EE", x"F2", x"EE", x"CD", x"A9", x"CD", x"D1", x"F1", x"F1", x"F1", x"F1", x"F1", x"D1", x"F1", x"A8", x"60", x"60", x"60", x"40", x"60", x"40", x"40", x"40", x"40", x"40", x"40", x"20", x"64", x"F1", x"CD", x"D2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"FB", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EA", x"EE", x"F2", x"F7", x"D7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"EA", x"C9", x"C9", x"CD", x"CD", x"CD", x"CD", x"CD", x"D6", x"FB", x"FA", x"DA", x"89", x"40", x"60", x"60", x"60", x"60", x"40", x"84", x"84", x"84", x"84", x"64", x"D1", x"D1", x"A8", x"AD", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"F1", x"F5", x"F5", x"F1", x"F1", x"DA", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EA", x"EE", x"F2", x"F3", x"F7", x"EE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"CD", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"64", x"40", x"40", x"40", x"60", x"AD", x"F2", x"F6", x"D1", x"AC", x"CD", x"F1", x"CD", x"AD", x"D6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F2", x"F1", x"F5", x"F1", x"F1", x"CD", x"CD", x"F1", x"F1", x"D1", x"CD", x"CD", x"FB", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"CE", x"EE", x"F2", x"F6", x"F7", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"C9", x"C9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"A9", x"CE", x"B2", x"D2", x"F7", x"F7", x"F7", x"D7", x"D2", x"D6", x"F6", x"D2", x"D6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F2", x"F2", x"F1", x"D1", x"D1", x"B1", x"D6", x"D6", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EE", x"EE", x"EE", x"F2", x"F7", x"EE", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F2", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"E9", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"FF", x"FF", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"F1", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"E9", x"F2", x"EE", x"F2", x"F7", x"EE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F2", x"EE", x"EE", x"EE", x"CD", x"AD", x"A9", x"85", x"C9", x"CD", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F2", x"FB", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F3", x"F7", x"F7", x"F2", x"F2", x"F2", x"F7", x"F7", x"F2", x"EE", x"EE", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EA", x"EE", x"EE", x"F2", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"C9", x"89", x"85", x"64", x"40", x"00", x"40", x"64", x"EE", x"EE", x"F2", x"FF", x"FB", x"FB", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F3", x"F7", x"F7", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"E9", x"F2", x"FB", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"EE", x"F2", x"F2", x"F7", x"EE", x"C9", x"65", x"44", x"20", x"00", x"00", x"65", x"89", x"89", x"CE", x"F2", x"F7", x"F2", x"CE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F3", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F6", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"89", x"20", x"20", x"00", x"40", x"A9", x"AD", x"A9", x"EE", x"F2", x"F2", x"F7", x"F7", x"F7", x"F2", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"85", x"00", x"00", x"20", x"A9", x"CE", x"F2", x"F7", x"F7", x"F6", x"F2", x"F7", x"F7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"85", x"20", x"40", x"A9", x"CE", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"EE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"85", x"EE", x"F7", x"F7", x"F2", x"F2", x"F3", x"F2", x"F7", x"F7", x"F7", x"F6", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"C9", x"EA", x"EE", x"EE", x"EE", x"EE", x"EE", x"F6", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"CE", x"F7", x"F7", x"F3", x"F6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"C9", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"EE", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F7", x"F2", x"EE", x"ED", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"EE", x"EE", x"F2", x"F7", x"F2", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"CE", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F3", x"F3", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"C5", x"C5", x"EE", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C5", x"EA", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"EE", x"C9", x"C9", x"CD", x"E9", x"C9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"EE", x"C9", x"C9", x"E9", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"ED", x"EE", x"C9", x"CA", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"C9", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CA", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"EE", x"EE", x"EA", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"EE", x"CD", x"ED", x"C9", x"CD", x"ED", x"ED", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"C5", x"E9", x"CD", x"CD", x"CD", x"CD", x"ED", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"C9", x"CD", x"D1", x"F1", x"CD", x"F1", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"CD", x"F1", x"F1", x"F1", x"F1", x"CD", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"CD", x"F1", x"F5", x"F5", x"F1", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"F5", x"F5", x"F5", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"F1", x"F5", x"F5", x"F5", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"F1", x"F1", x"F5", x"F5", x"F5", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F1", x"F1", x"F1", x"F1", x"F5", x"F1", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"F1", x"CD", x"CD", x"CD", x"CD", x"AC", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F1", x"F1", x"ED", x"AD", x"AD", x"AC", x"CD", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"CD", x"F1", x"F1", x"ED", x"CD", x"AD", x"CD", x"CD", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"CD", x"AD", x"F1", x"F1", x"F1", x"D1", x"CD", x"F1", x"F1", x"ED", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"CD", x"CD", x"CC", x"CD", x"CD", x"CD", x"CC", x"CD", x"CD", x"CD", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B1", x"D6", x"D6", x"D6", x"B1", x"B1", x"D2", x"D1", x"B1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
);
constant PinkKick_bmp: PinkKick_bmp_array := (
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000011110000000000000000000000000000000000000000000000000000000000000000000000000"),
("000001111111110000000001111111100000000000000000000000000000000000000000000000000000"),
("000111111111111100000111111111110000000000000000000000000000000000000000000000000000"),
("000010111111111100001111111111111000000000000000000000000000000000000000000000000000"),
("000011111111111111111111111111111000111110000000000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111100000000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111000000000000000000000000000000000000000"),
("001111101111000001111111111111111111111111111100000000000000000000000000000000000000"),
("001110001000000011111111111111111111111111111110000000000000000000000000000000000000"),
("001100010000101111111111111111111111111111111110000000000000000000000000000001110000"),
("001100010011111111111111111111111111111111111100000000000000000000000000000011110000"),
("000100010011111111111111111111111111111110000000000000000000000000000000000011110000"),
("000100000011111111111111111111111111111100000000000000000000000000000000000111111000"),
("000010000111111111111111111111111111111100000000000000000000000000000000001111111000"),
("000000000111111111111111111111111111111111000000000000000000000000000000001111111000"),
("000000000111111111111111111111111111111111111111111111111110000000000000011111111000"),
("000000001111111111111111111111111111111111111111111111111110000000000000111111110000"),
("000000001111111111111111111111111111111111111111111111111111000000000001111111110000"),
("000000001111111111111111111111111111111111111111111111111111100000000011111111110000"),
("000000001111111111111111111111111111111111111111111111111111101111111111111111111000"),
("000000001111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000000000111111111111111111111111111110000000111111111111111111111111111111111111100"),
("000000000011111111111111111111111111000000000111111111111111111111111111111111100000"),
("000000000001111111111111111111111111000000010011111111111111111111111111100000000000"),
("000000000000111111111111111111111110000011111111111111111111111111111111100000000000"),
("000000000000011111111111111111111110111111111111111111111111111111111111100000000000"),
("000000000000001111111111111111111111111111111111111111111111111111111000000000000000"),
("000000000000000111111111111111111111111111111111111111111111111111000000000000000000"),
("000000000000000011111111111111111111111111111111111111111111111000000000000000000000"),
("000000000000000001111111111111111111111111111111111111111111100000000000000000000000"),
("000000000000000001111111111111111111111111111111111111111111000000000000000000000000"),
("000000000000000001111111111111111111111111111111111111111000000000000000000000000000"),
("000000000000000000111111111111111111111111111111100000000000000000000000000000000000"),
("000000000000000000111111111111111111111111111110000000000000000000000000000000000000"),
("000000000000000000111111111111111111111111111000000000000000000000000000000000000000"),
("000000000000000001111111111111111111111111100000000000000000000000000000000000000000"),
("000000000000000001111111111111111111111111000000000000000000000000000000000000000000"),
("000000000000000001111111111111111111111000000000000000000000000000000000000000000000"),
("000000000000000000111111111111111111100000000000000000000000000000000000000000000000"),
("000000000000000000111111111111111111000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111111110000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111111110000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111111110000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111111100000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111111100000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111111000000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111111000000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111111000000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111110000000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111110000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111110000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111100000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111100000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111100000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111100000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111100000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111100000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111100000000000000000000000000000000000000000000000000000"),
("000000000000000001111111111111000000000000000000000000000000000000000000000000000000"),
("000000000000000001111111111111000000000000000000000000000000000000000000000000000000"),
("000000000000000001111111111111000000000000000000000000000000000000000000000000000000"),
("000000000000000001111111111110000000000000000000000000000000000000000000000000000000"),
("000000000000000001111111111110000000000000000000000000000000000000000000000000000000"),
("000000000000000011111111111110000000000000000000000000000000000000000000000000000000"),
("000000000000000011111111111100000000000000000000000000000000000000000000000000000000"),
("000000000000000011111111110000000000000000000000000000000000000000000000000000000000"),
("000000000000000011111111110000000000000000000000000000000000000000000000000000000000"),
("000000000000000000011111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000000011111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000000011111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000000011111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000000111111110000000000000000000000000000000000000000000000000000000000"),
("000000000000000000111111110000000000000000000000000000000000000000000000000000000000"),
("000000000000000001111111110000000000000000000000000000000000000000000000000000000000"),
("000000000000000011111111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000111111111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000111111111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000011111111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);
constant PinkDucking_X_size : integer := 91;
constant PinkDucking_Y_size : integer := 83;
type PinkDucking_color_array is array(0 to PinkDucking_Y_size - 1 , 0 to PinkDucking_X_size - 1) of std_logic_vector(7 downto 0);
type PinkDucking_bmp_array is array(0 to PinkDucking_Y_size - 1 , 0 to PinkDucking_X_size - 1) of std_logic;
constant PinkDucking_colors: PinkDucking_color_array := (
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"D6", x"D6", x"D6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D2", x"AD", x"88", x"84", x"64", x"84", x"84", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"A9", x"64", x"84", x"88", x"88", x"88", x"88", x"88", x"84", x"84", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"88", x"68", x"88", x"84", x"88", x"84", x"64", x"CC", x"CC", x"88", x"88", x"64", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"88", x"88", x"88", x"A8", x"CD", x"88", x"88", x"64", x"68", x"68", x"D1", x"D1", x"88", x"84", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"FB", x"FB", x"FB", x"DA", x"B1", x"84", x"A8", x"88", x"84", x"D1", x"F5", x"A8", x"D1", x"D1", x"68", x"00", x"F6", x"FA", x"CD", x"64", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"FB", x"F7", x"FB", x"FF", x"FB", x"F2", x"F2", x"EE", x"EE", x"C9", x"C9", x"C9", x"A8", x"CC", x"CD", x"CC", x"A8", x"D1", x"D1", x"D1", x"F6", x"F6", x"AD", x"24", x"89", x"F1", x"AD", x"92", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F7", x"F7", x"F2", x"F2", x"EE", x"CE", x"CA", x"CE", x"F2", x"CD", x"C9", x"C9", x"A8", x"CD", x"F1", x"F1", x"F1", x"F1", x"CD", x"CD", x"F5", x"FA", x"FA", x"FA", x"F5", x"CD", x"D1", x"CD", x"CD", x"DB", x"D6", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F2", x"CD", x"F2", x"F7", x"F2", x"F7", x"F6", x"EE", x"EE", x"F7", x"F2", x"CD", x"CD", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"CD", x"D1", x"FA", x"FA", x"F6", x"FA", x"F6", x"F1", x"D5", x"D1", x"EE", x"CD", x"C9", x"FB", x"FB", x"F7", x"F7", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F5", x"F6", x"D2", x"D2", x"F2", x"F2", x"F7", x"F2", x"EE", x"F2", x"F7", x"D2", x"CD", x"F1", x"D1", x"F5", x"F5", x"F1", x"F1", x"F6", x"D1", x"CD", x"CD", x"F5", x"F6", x"F6", x"FA", x"D5", x"A8", x"AD", x"CD", x"F6", x"F2", x"F6", x"F2", x"EE", x"EE", x"EE", x"C9", x"CD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"FA", x"FA", x"F2", x"F2", x"F2", x"F7", x"F7", x"D2", x"EE", x"F7", x"F7", x"F2", x"64", x"88", x"F1", x"F1", x"F1", x"F5", x"F6", x"F1", x"F1", x"F1", x"ED", x"AC", x"CD", x"F5", x"D1", x"D1", x"AD", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F2", x"EE", x"CD", x"CD", x"C5", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F1", x"F6", x"F6", x"F2", x"F2", x"F2", x"D7", x"F7", x"F2", x"EE", x"F7", x"F7", x"F2", x"60", x"00", x"6D", x"D1", x"D1", x"F5", x"CD", x"D1", x"F1", x"D1", x"88", x"64", x"44", x"CD", x"CE", x"CD", x"CE", x"F7", x"F7", x"F7", x"F7", x"F6", x"F3", x"F2", x"F2", x"F2", x"F5", x"D1", x"C9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"D1", x"F5", x"D1", x"D2", x"F3", x"F2", x"F7", x"F7", x"D2", x"EE", x"F7", x"F7", x"D2", x"60", x"00", x"00", x"24", x"44", x"24", x"20", x"24", x"24", x"24", x"00", x"00", x"20", x"C9", x"F7", x"EE", x"EE", x"F7", x"F7", x"D7", x"D7", x"F7", x"F2", x"F2", x"F1", x"FA", x"FA", x"FA", x"ED", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F1", x"D1", x"F1", x"F2", x"F2", x"F7", x"D7", x"F2", x"EE", x"F7", x"F7", x"F2", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"CE", x"F7", x"F2", x"EE", x"F7", x"F2", x"F7", x"F7", x"F6", x"F2", x"F5", x"F1", x"F6", x"F1", x"F1", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"F1", x"F1", x"F2", x"F2", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F2", x"64", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"EE", x"F7", x"F2", x"EE", x"F7", x"EE", x"F2", x"F7", x"F2", x"ED", x"F1", x"F5", x"F6", x"F1", x"CD", x"CD", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F5", x"F1", x"F2", x"F2", x"F2", x"F7", x"F2", x"EE", x"F7", x"F7", x"F7", x"69", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"A9", x"D7", x"F7", x"EE", x"F2", x"D7", x"F2", x"F2", x"F2", x"CD", x"CD", x"F6", x"FA", x"FA", x"FA", x"F6", x"D1", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"ED", x"EE", x"F2", x"F2", x"F7", x"F7", x"EE", x"F2", x"F7", x"F7", x"AE", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"44", x"69", x"F3", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"EE", x"EE", x"CD", x"CD", x"F1", x"F9", x"FA", x"FA", x"FA", x"FA", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"F1", x"F1", x"ED", x"EE", x"F2", x"F2", x"F7", x"F2", x"EE", x"F7", x"F7", x"F7", x"65", x"00", x"00", x"00", x"00", x"20", x"44", x"65", x"AE", x"D2", x"F7", x"F7", x"F2", x"F2", x"F7", x"D7", x"F7", x"F3", x"F2", x"EE", x"AD", x"AD", x"CD", x"F1", x"F6", x"FA", x"F6", x"FA", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"D6", x"D6", x"A8", x"AC", x"ED", x"CD", x"CD", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F7", x"F7", x"D2", x"69", x"00", x"00", x"44", x"CE", x"F2", x"F7", x"F7", x"F7", x"F2", x"EE", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"CD", x"CD", x"A8", x"A8", x"AD", x"ED", x"F6", x"FA", x"FA", x"FA", x"F1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"D1", x"A8", x"84", x"A8", x"A8", x"A8", x"C9", x"EE", x"EE", x"F2", x"F2", x"EE", x"CE", x"F2", x"F7", x"F7", x"89", x"65", x"EE", x"F7", x"F7", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F1", x"F1", x"D1", x"CD", x"AD", x"AC", x"CD", x"F1", x"F5", x"F5", x"F1", x"CD", x"D1", x"FA", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D6", x"F6", x"D5", x"F6", x"F6", x"D6", x"FB", x"DA", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AC", x"D1", x"CD", x"D1", x"CD", x"A8", x"AD", x"A8", x"AD", x"84", x"A9", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F7", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"EE", x"C9", x"CD", x"F1", x"D1", x"CD", x"CD", x"CD", x"CD", x"CD", x"F1", x"F5", x"D1", x"D1", x"F5", x"F6", x"F6", x"FB", x"FB", x"FB", x"DB", x"DA", x"DB", x"DB", x"DB", x"DB", x"D6", x"D5", x"F5", x"F1", x"A8", x"A8", x"AD", x"44", x"D1", x"AD", x"FB", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F6", x"CD", x"D1", x"D1", x"D1", x"F5", x"AD", x"F5", x"D1", x"C9", x"F2", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"ED", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"E9", x"D1", x"AD", x"CC", x"CD", x"A9", x"CD", x"D1", x"CD", x"AC", x"CD", x"F5", x"F5", x"F1", x"F1", x"F5", x"F5", x"F5", x"D5", x"D1", x"CD", x"88", x"64", x"64", x"64", x"64", x"B1", x"FA", x"FA", x"D1", x"44", x"69", x"B1", x"6D", x"D1", x"88", x"FB", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"68", x"D1", x"F1", x"CD", x"F5", x"F5", x"F1", x"F1", x"F5", x"CD", x"A9", x"E9", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"C9", x"C9", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"CE", x"EE", x"EE", x"EE", x"D7", x"FF", x"FB", x"DA", x"AD", x"A8", x"CD", x"CD", x"D5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"64", x"40", x"40", x"40", x"40", x"AD", x"F1", x"F1", x"AD", x"44", x"8D", x"D5", x"F1", x"AD", x"B1", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"69", x"84", x"A8", x"A8", x"A8", x"AD", x"AD", x"AD", x"A8", x"60", x"20", x"40", x"85", x"CE", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"E9", x"EE", x"EE", x"EE", x"EE", x"EA", x"EE", x"EE", x"EE", x"E9", x"C9", x"EE", x"F2", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"CD", x"CD", x"F5", x"F6", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"88", x"60", x"60", x"40", x"40", x"AD", x"F1", x"D1", x"CD", x"44", x"AD", x"F5", x"F5", x"AD", x"DA", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"88", x"89", x"88", x"84", x"84", x"60", x"84", x"84", x"60", x"00", x"00", x"24", x"65", x"A9", x"C9", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"E9", x"EE", x"EE", x"A9", x"A5", x"A5", x"A9", x"CE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"AC", x"CD", x"F1", x"F5", x"F5", x"F6", x"F6", x"F6", x"F6", x"F5", x"F5", x"F5", x"F5", x"F5", x"64", x"40", x"40", x"40", x"40", x"88", x"D5", x"F6", x"F5", x"68", x"68", x"F1", x"D1", x"AD", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F6", x"F2", x"ED", x"C9", x"EE", x"EE", x"A9", x"64", x"60", x"00", x"00", x"00", x"20", x"60", x"64", x"85", x"85", x"69", x"89", x"64", x"60", x"64", x"40", x"20", x"64", x"89", x"D2", x"FB", x"FB", x"FB", x"FB", x"F7", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D6", x"FA", x"D6", x"F1", x"D5", x"D5", x"F1", x"D1", x"D1", x"D1", x"CD", x"CD", x"A8", x"64", x"40", x"20", x"20", x"20", x"40", x"84", x"A8", x"C9", x"44", x"00", x"84", x"A8", x"B1", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F2", x"F7", x"F2", x"EE", x"E9", x"E9", x"C9", x"85", x"44", x"24", x"20", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"44", x"A5", x"A5", x"EA", x"EE", x"CE", x"EE", x"F2", x"F3", x"F2", x"D2", x"EE", x"FB", x"FB", x"FB", x"F7", x"F6", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"D6", x"FB", x"FB", x"FB", x"FB", x"DA", x"DA", x"DA", x"AD", x"89", x"89", x"89", x"D6", x"8D", x"68", x"89", x"69", x"69", x"89", x"8D", x"FB", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"F7", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F3", x"D2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"20", x"00", x"00", x"00", x"00", x"A5", x"EE", x"EA", x"EA", x"EE", x"EE", x"F2", x"F7", x"EE", x"EE", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"F7", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"F7", x"F7", x"F7", x"F3", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"CE", x"44", x"00", x"00", x"45", x"65", x"20", x"44", x"CE", x"EE", x"E9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F6", x"F7", x"F7", x"D7", x"F7", x"D7", x"F3", x"F6", x"F7", x"D7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"EE", x"EA", x"EE", x"CD", x"EE", x"EE", x"65", x"00", x"20", x"A9", x"F2", x"EE", x"20", x"00", x"44", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"D7", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F3", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F2", x"F2", x"EE", x"EE", x"89", x"00", x"20", x"65", x"EE", x"EE", x"EE", x"65", x"00", x"00", x"89", x"E9", x"E9", x"EE", x"EE", x"F2", x"F7", x"F3", x"F3", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F2", x"F2", x"F7", x"F7", x"D7", x"D7", x"F7", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"F2", x"F3", x"F7", x"F7", x"F7", x"F3", x"D7", x"F7", x"F7", x"F3", x"F7", x"D7", x"F3", x"F2", x"F2", x"F2", x"F6", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"89", x"00", x"00", x"A5", x"C9", x"E9", x"C9", x"C9", x"20", x"20", x"85", x"CE", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"F2", x"F2", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F3", x"EE", x"EE", x"F7", x"F7", x"F7", x"D7", x"F7", x"F2", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"EE", x"F2", x"F2", x"F7", x"D7", x"EE", x"F6", x"F7", x"F2", x"F2", x"F2", x"F7", x"EE", x"EE", x"F2", x"F6", x"D7", x"F2", x"F2", x"EE", x"ED", x"ED", x"EE", x"EE", x"85", x"00", x"20", x"C9", x"C9", x"C9", x"EE", x"C9", x"20", x"00", x"44", x"A9", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"EE", x"F2", x"F2", x"F7", x"F2", x"F2", x"F2", x"F7", x"F7", x"F2", x"F2", x"F2", x"CE", x"ED", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"20", x"00", x"85", x"EE", x"EE", x"EE", x"EE", x"EE", x"A9", x"00", x"00", x"89", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"F2", x"F6", x"F3", x"D7", x"F7", x"D7", x"F2", x"F2", x"EE", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F7", x"F7", x"F3", x"F2", x"CE", x"C9", x"C9", x"EE", x"EE", x"EE", x"EE", x"EE", x"E9", x"E9", x"A5", x"00", x"00", x"A5", x"E9", x"C5", x"C5", x"C9", x"C9", x"C5", x"00", x"00", x"89", x"EE", x"EA", x"ED", x"EA", x"EE", x"EE", x"EE", x"EE", x"C9", x"C5", x"C9", x"EA", x"EA", x"EE", x"EA", x"C9", x"EE", x"EE", x"F2", x"F3", x"F7", x"D7", x"F7", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"F7", x"F7", x"F7", x"F2", x"C9", x"C9", x"E9", x"C9", x"C9", x"EE", x"EE", x"F2", x"D2", x"A9", x"00", x"00", x"A9", x"CE", x"CE", x"CE", x"CE", x"CE", x"AD", x"00", x"00", x"89", x"EE", x"CE", x"CE", x"CE", x"D2", x"CE", x"F2", x"F2", x"D2", x"CE", x"D2", x"F2", x"F2", x"D2", x"C9", x"C5", x"E9", x"EE", x"F2", x"F7", x"F7", x"D7", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"E9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"CE", x"F2", x"F2", x"C9", x"EE", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"DB", x"24", x"24", x"D7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"24", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"C5", x"EE", x"D2", x"F7", x"D7", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F7", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"E9", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"D7", x"F7", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"EE", x"F2", x"F7", x"F7", x"F2", x"ED", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"E9", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F6", x"F7", x"CE", x"EE", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EE", x"CD", x"CD", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"EA", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"EE", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"CD", x"EE", x"CE", x"F7", x"EE", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F6", x"D1", x"CD", x"ED", x"ED", x"ED", x"ED", x"CD", x"ED", x"EE", x"EE", x"EE", x"F6", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"CD", x"CE", x"F2", x"E9", x"C9", x"CD", x"EA", x"CD", x"ED", x"CD", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"ED", x"F1", x"F1", x"F1", x"F1", x"CD", x"D6", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"D2", x"CD", x"ED", x"CD", x"CD", x"CD", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"F1", x"F5", x"F1", x"F1", x"ED", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"F1", x"F1", x"F1", x"F1", x"CD", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"F1", x"F5", x"F5", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AD", x"F1", x"F1", x"F1", x"F5", x"F1", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"F1", x"F5", x"F5", x"F1", x"F1", x"F1", x"D1", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F5", x"F1", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"D1", x"F1", x"F5", x"F5", x"F1", x"F1", x"F1", x"F1", x"F1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F1", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"F5", x"F1", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F1", x"F5", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"F1", x"F1", x"F1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FB", x"DB", x"FB", x"D6", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"D1", x"D1", x"D2", x"D5", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"D1", x"D1", x"ED", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"D6", x"FB", x"FB", x"FB", x"DB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FB", x"D2", x"CD", x"D1", x"F5", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"ED", x"CD", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"F5", x"F1", x"F5", x"F1", x"F1", x"F1", x"D1", x"D1", x"CD", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FB", x"CC", x"84", x"CD", x"D1", x"CD", x"CC", x"D1", x"D1", x"D1", x"CD", x"D2", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F5", x"F5", x"F5", x"F6", x"D6", x"F1", x"D1", x"F6", x"D5", x"D1", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FB", x"DA", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
);
constant PinkDucking_bmp: PinkDucking_bmp_array := (
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000"),
("0000000000000000000000000000000000111111111111111111111100000000000000000000000000000000000"),
("0000000000000000000000000101110111111111111111111111111110000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111111111110000000000000000000000000000000000"),
("0000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000"),
("0000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000"),
("0000000000000000000011111111111111111111111111111111111111111111000000000000000000000000000"),
("0000000000000000000011111111111111111111111111111111111111111111000000000000000000000000000"),
("0000000000000000000011111111111111111111111111111111111111111111000000000000000000000000000"),
("0000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000"),
("0000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000"),
("0000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000"),
("0000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000"),
("0000000000000000000000111111111111111111111111111111111111111111100000000000000000000000000"),
("0000000000000000000111111111111111111111111111111111111111111111110000000000000000000000000"),
("0000000000000000001111111111111111111111111111111111111111111111111110000000000011111111100"),
("0000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110"),
("0000000000000000011111111111111111111111111111111111111111111111111111111111111111111111110"),
("0000000000000000011111111111111111111111111111111111110111111111111111111111111111111111100"),
("0000000000000000011111111111111111111111111111111111100000111111111111111111111111111111100"),
("0000000000000000000111111111111111111111111111111100000000011111111111111111111111111111000"),
("0000000000000000000001111111111111111111111111111111111000001111111111111111111111111111000"),
("0000000000000000111111111111111111111111111111111111111111110000111111111111111111111111000"),
("0000000000000111111111111111111111111111111111111111111111111111111110000000000000100000000"),
("0000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("0000000011111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("0000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000"),
("0000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000"),
("0000000111111111111111111111111111111111111111111111111111111111111111111000000000000000000"),
("0000000111111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("0000000011111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("0000000011111111111111111111111111111111111111111111111111111111111111111110000000000000000"),
("0000000011111111111111111111100011110000011110000000000000111111111111111110000000000000000"),
("0000000011111111111111110000000000100000001100000000000000111111111111111111000000000000000"),
("0000000011111111111111110000000000000000000000000000000000011111111111111111100000000000000"),
("0000000011111111111111100000000000000000000000000000000000011111111111111111110000000000000"),
("0000000011111111111111100000000000000000000000000000000000001111111111111111100000000000000"),
("0000000011111111111111100000000000000000000000000000000000000111111111111000000000000000000"),
("0000000000111111111110000000000000000000000000000000000000000011111111110000000000000000000"),
("0000000000111111110000000000000000000000000000000000000000000000111111110000000000000000000"),
("0000000000111111100000000000000000000000000000000000000000000001111111100000000000000000000"),
("0000000001111111110000000000000000000000000000000000000000000111111111100000000000000000000"),
("0000000011111111111000000000000000000000000000000000000000001111111111100000000000000000000"),
("0000000111111111111100000000000000000000000000000000000000001111111111110000000000000000000"),
("0000000111111111111100000000000000000000000000000000000000001111111111110000000000000000000"),
("0001111111111111111000000000000000000000000000000000000000000111111111111111110000000000000"),
("0111111111111111000000000000000000000000000000000000000000000000011111111111111000000000000"),
("0111111111111100000000000000000000000000000000000000000000000000001111111111111000000000000"),
("0011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000")
);
constant PinkHitted_X_size : integer := 63;
constant PinkHitted_Y_size : integer := 83;
type PinkHitted_color_array is array(0 to PinkHitted_Y_size - 1 , 0 to PinkHitted_X_size - 1) of std_logic_vector(7 downto 0);
type PinkHitted_bmp_array is array(0 to PinkHitted_Y_size - 1 , 0 to PinkHitted_X_size - 1) of std_logic;
constant PinkHitted_colors: PinkHitted_color_array := (
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AD", x"84", x"88", x"84", x"88", x"84", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"84", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"D6", x"88", x"A8", x"AD", x"AC", x"88", x"88", x"88", x"84", x"88", x"88", x"84", x"B1", x"FF", x"FF", x"FF", x"FF", x"DA", x"FF", x"AD", x"8D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"8D", x"88", x"AC", x"F5", x"B1", x"CC", x"D1", x"88", x"88", x"8C", x"88", x"84", x"84", x"D6", x"FF", x"FF", x"FF", x"D6", x"B1", x"B1", x"88", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FA", x"88", x"88", x"B1", x"49", x"D1", x"F6", x"F5", x"88", x"D1", x"FA", x"F1", x"88", x"84", x"AD", x"FB", x"DB", x"DA", x"A8", x"88", x"88", x"DA", x"D6", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"B2", x"88", x"A8", x"B1", x"00", x"8D", x"FA", x"F6", x"AC", x"AC", x"F6", x"F5", x"A8", x"A8", x"A4", x"A8", x"8C", x"A8", x"84", x"88", x"AD", x"B1", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"DB", x"B1", x"88", x"A8", x"D1", x"B1", x"44", x"D1", x"F5", x"F6", x"F6", x"AC", x"CC", x"F1", x"CD", x"F1", x"A8", x"A4", x"A8", x"A8", x"88", x"88", x"AD", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F6", x"F1", x"CD", x"F1", x"FA", x"F6", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"B1", x"D6", x"D6", x"D6", x"6D", x"AD", x"68", x"F1", x"F1", x"F6", x"FA", x"F5", x"F1", x"F5", x"CD", x"F5", x"F5", x"CD", x"84", x"84", x"88", x"88", x"88", x"88", x"B1", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"CD", x"A8", x"D1", x"F1", x"F1", x"AD", x"CD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"AD", x"FF", x"FF", x"FF", x"DA", x"A8", x"CD", x"F1", x"F6", x"FA", x"FA", x"FA", x"F6", x"F6", x"F1", x"F1", x"F6", x"F5", x"D1", x"C9", x"CD", x"D2", x"D2", x"D2", x"D2", x"F7", x"F2", x"EE", x"F6", x"FB", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"AD", x"F1", x"A8", x"D1", x"F6", x"D1", x"CD", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F5", x"F1", x"F1", x"F6", x"F1", x"F5", x"FA", x"F5", x"D1", x"F5", x"F1", x"F5", x"FA", x"F5", x"CD", x"C9", x"C9", x"A5", x"A5", x"F2", x"F7", x"F2", x"EE", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"F5", x"FB", x"92", x"44", x"AD", x"A8", x"AD", x"F5", x"CD", x"CD", x"CD", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F6", x"D1", x"D1", x"FB", x"F6", x"F5", x"F6", x"F1", x"AD", x"F5", x"F5", x"F6", x"F6", x"FA", x"F6", x"F1", x"F1", x"88", x"48", x"A5", x"C9", x"EE", x"F2", x"F2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F5", x"F1", x"44", x"00", x"44", x"88", x"CD", x"AC", x"88", x"CD", x"F1", x"CD", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"CC", x"D1", x"F1", x"F6", x"D5", x"CD", x"D1", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"F1", x"F1", x"CD", x"88", x"20", x"A5", x"EE", x"F2", x"CE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F1", x"D1", x"44", x"00", x"00", x"64", x"A8", x"CD", x"CD", x"AD", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"ED", x"AD", x"CD", x"CD", x"CD", x"D2", x"F7", x"F6", x"F6", x"F6", x"F2", x"ED", x"F6", x"F5", x"CD", x"CD", x"AD", x"24", x"00", x"20", x"A5", x"EE", x"F2", x"EE", x"CA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"F5", x"D1", x"44", x"00", x"00", x"44", x"44", x"68", x"AC", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"C9", x"E9", x"EE", x"EE", x"F2", x"F6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"F1", x"D1", x"44", x"00", x"00", x"00", x"24", x"A5", x"EE", x"F2", x"C9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"8C", x"CD", x"F1", x"F1", x"AD", x"AD", x"89", x"20", x"00", x"00", x"44", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"FB", x"F2", x"C9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F3", x"F7", x"F7", x"F7", x"F2", x"F2", x"AE", x"44", x"20", x"00", x"00", x"20", x"A5", x"EE", x"F2", x"F7", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FB", x"B1", x"40", x"40", x"84", x"A8", x"CC", x"D1", x"F1", x"CD", x"64", x"44", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"F7", x"F6", x"EE", x"CD", x"8D", x"CE", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F7", x"F7", x"F6", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F2", x"A9", x"44", x"00", x"00", x"44", x"E9", x"F3", x"CD", x"CD", x"F6", x"FB", x"FF", x"FF", x"D6", x"CD", x"A8", x"40", x"20", x"40", x"40", x"64", x"A8", x"C8", x"AC", x"8C", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"F6", x"F2", x"CE", x"C9", x"64", x"24", x"00", x"40", x"69", x"69", x"8D", x"F2", x"F6", x"F3", x"F3", x"D7", x"F7", x"D7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F3", x"F7", x"F7", x"F2", x"89", x"00", x"20", x"A5", x"D2", x"F2", x"C9", x"F1", x"CD", x"C9", x"CD", x"F1", x"F5", x"AC", x"40", x"20", x"40", x"40", x"20", x"40", x"40", x"60", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"F6", x"E9", x"C9", x"44", x"24", x"D1", x"D1", x"B1", x"91", x"00", x"69", x"F3", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F2", x"F3", x"F7", x"F2", x"89", x"00", x"20", x"A9", x"F2", x"EE", x"CD", x"CD", x"CD", x"F1", x"F5", x"F5", x"F1", x"88", x"64", x"40", x"40", x"20", x"40", x"40", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"F6", x"C9", x"68", x"B1", x"D6", x"FA", x"FA", x"FA", x"FA", x"D5", x"F6", x"8D", x"44", x"AE", x"D7", x"D7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"89", x"00", x"85", x"F2", x"EE", x"C9", x"CD", x"F1", x"F1", x"F1", x"F1", x"F5", x"F1", x"CC", x"84", x"84", x"64", x"88", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"EE", x"64", x"B1", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F1", x"D1", x"68", x"EE", x"F7", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F3", x"EE", x"F2", x"F6", x"F7", x"89", x"A5", x"EE", x"EE", x"C9", x"ED", x"F1", x"F1", x"ED", x"D1", x"ED", x"F1", x"D1", x"F1", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"EE", x"44", x"B1", x"F5", x"F5", x"FA", x"F6", x"FA", x"F6", x"F1", x"F1", x"F6", x"FA", x"FA", x"F1", x"EE", x"F2", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"F2", x"F7", x"F7", x"CE", x"EE", x"EE", x"E9", x"EE", x"C9", x"CD", x"CD", x"CD", x"CD", x"ED", x"F1", x"ED", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"F2", x"44", x"B1", x"F5", x"F1", x"F5", x"F5", x"F6", x"F5", x"F1", x"F1", x"F6", x"FA", x"FA", x"F6", x"F1", x"EE", x"F2", x"EE", x"F3", x"D7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F3", x"EE", x"EE", x"F7", x"F2", x"C9", x"CE", x"E9", x"F2", x"C9", x"A9", x"CD", x"D1", x"ED", x"ED", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"F2", x"C9", x"CD", x"F1", x"F1", x"F1", x"F1", x"F1", x"F5", x"F6", x"F6", x"F6", x"F6", x"FA", x"FA", x"F5", x"CD", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"F2", x"EE", x"C9", x"C9", x"EE", x"C5", x"CD", x"D1", x"ED", x"D1", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"F2", x"C9", x"CD", x"ED", x"F1", x"F1", x"F1", x"F6", x"FA", x"FA", x"F6", x"F5", x"F1", x"F6", x"F5", x"CD", x"CD", x"CE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"CE", x"C9", x"CE", x"CE", x"A5", x"C5", x"C9", x"A4", x"AC", x"AD", x"AD", x"AC", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"CD", x"F5", x"F5", x"F6", x"F5", x"F6", x"F6", x"F6", x"F6", x"F1", x"F1", x"F1", x"F1", x"F1", x"CD", x"CD", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"CE", x"C9", x"A9", x"80", x"40", x"40", x"40", x"40", x"20", x"84", x"CD", x"F1", x"CD", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"F5", x"F6", x"F5", x"F1", x"F1", x"F1", x"F5", x"F5", x"F5", x"FA", x"F6", x"FA", x"F6", x"F5", x"F5", x"ED", x"CD", x"CD", x"A9", x"89", x"60", x"40", x"40", x"40", x"40", x"60", x"40", x"40", x"40", x"D1", x"F6", x"F5", x"D1", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F5", x"F5", x"F5", x"F1", x"CD", x"F5", x"FA", x"FA", x"FA", x"F6", x"FA", x"F6", x"F6", x"F6", x"F6", x"D1", x"AD", x"40", x"40", x"60", x"40", x"40", x"40", x"60", x"60", x"60", x"40", x"AD", x"F6", x"F5", x"F6", x"F1", x"D1", x"D1", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"F1", x"F6", x"F5", x"CD", x"CD", x"F5", x"F5", x"F5", x"F6", x"F5", x"F6", x"F6", x"F6", x"FA", x"F6", x"64", x"40", x"60", x"40", x"40", x"60", x"60", x"40", x"40", x"40", x"64", x"F6", x"F5", x"F1", x"F6", x"F5", x"F1", x"CD", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"A9", x"CD", x"F5", x"F5", x"CD", x"CD", x"F1", x"F5", x"FA", x"F6", x"FA", x"F6", x"FA", x"FA", x"F6", x"40", x"60", x"60", x"40", x"40", x"60", x"40", x"60", x"60", x"40", x"64", x"F6", x"F6", x"F6", x"F1", x"F1", x"D1", x"F6", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C5", x"A9", x"CD", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F6", x"F6", x"FA", x"F6", x"F6", x"F6", x"40", x"40", x"60", x"40", x"40", x"40", x"40", x"40", x"40", x"64", x"F5", x"F6", x"F1", x"F5", x"F5", x"F5", x"D1", x"AD", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C5", x"C5", x"CD", x"F5", x"F1", x"F1", x"F1", x"F1", x"F1", x"F5", x"F5", x"F1", x"F5", x"F1", x"88", x"40", x"60", x"60", x"40", x"40", x"40", x"44", x"20", x"CD", x"D1", x"D1", x"F5", x"F6", x"CD", x"CD", x"D1", x"D1", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"D6", x"CD", x"F1", x"F5", x"F5", x"F1", x"F1", x"F1", x"F1", x"F5", x"F5", x"F1", x"D1", x"CD", x"84", x"64", x"40", x"40", x"20", x"64", x"A9", x"84", x"44", x"44", x"24", x"8D", x"F5", x"D1", x"C9", x"CD", x"CE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"CD", x"CD", x"D1", x"F1", x"F1", x"CD", x"CD", x"CD", x"CD", x"CD", x"CD", x"CD", x"CD", x"CE", x"CD", x"CD", x"EE", x"ED", x"A9", x"00", x"00", x"20", x"44", x"AD", x"CD", x"F2", x"F2", x"EE", x"C9", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"CD", x"CD", x"CD", x"AD", x"C9", x"CD", x"F2", x"F3", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"CD", x"00", x"00", x"64", x"40", x"20", x"A9", x"EE", x"EE", x"C9", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"C9", x"EE", x"C9", x"CD", x"ED", x"EE", x"EA", x"EE", x"F7", x"D7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"CD", x"00", x"00", x"65", x"64", x"00", x"24", x"C9", x"EE", x"ED", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"CE", x"C9", x"EA", x"EA", x"EE", x"F2", x"EE", x"E9", x"EE", x"F3", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"EE", x"C9", x"44", x"00", x"00", x"84", x"20", x"00", x"20", x"CE", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"ED", x"E9", x"C9", x"EE", x"F2", x"F2", x"F2", x"EE", x"C9", x"ED", x"CE", x"CE", x"CE", x"E9", x"C9", x"C9", x"C9", x"E9", x"A9", x"00", x"00", x"44", x"64", x"00", x"00", x"44", x"CE", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"C9", x"C9", x"E9", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"64", x"00", x"00", x"A9", x"89", x"00", x"00", x"24", x"CE", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"C9", x"CD", x"EE", x"EE", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"E9", x"85", x"00", x"00", x"24", x"AE", x"20", x"00", x"00", x"24", x"F2", x"F2", x"ED", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"E9", x"E9", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"F2", x"EE", x"C9", x"C9", x"E9", x"65", x"00", x"00", x"AE", x"AE", x"20", x"00", x"44", x"F7", x"D7", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"C5", x"EE", x"F2", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F2", x"E9", x"C9", x"EE", x"EE", x"65", x"00", x"00", x"24", x"F7", x"B2", x"69", x"CE", x"D7", x"F7", x"F3", x"F2", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"E9", x"EE", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"E9", x"C9", x"EE", x"EE", x"65", x"00", x"20", x"AD", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"F2", x"EE", x"F7", x"D7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"E9", x"ED", x"EE", x"EE", x"C9", x"44", x"A9", x"F2", x"D7", x"D7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"C9", x"EE", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"C9", x"E9", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"D7", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F2", x"C9", x"C9", x"EE", x"EE", x"F2", x"F2", x"F6", x"F7", x"F2", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"E9", x"EE", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"C9", x"CE", x"EA", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F2", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"F2", x"C9", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F7", x"D7", x"F2", x"F2", x"F7", x"D7", x"F7", x"F7", x"D7", x"F7", x"F7", x"D7", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E9", x"F2", x"F2", x"D7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F3", x"F2", x"C9", x"FF", x"FF", x"EE", x"EE", x"F2", x"EE", x"F2", x"F7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"EE", x"F2", x"F7", x"D7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"C9", x"FF", x"FF", x"FB", x"E9", x"EE", x"F2", x"F2", x"F7", x"F7", x"F3", x"F7", x"D7", x"F7", x"D7", x"F7", x"F2", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"E9", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"EE", x"C5", x"FF", x"FF", x"FF", x"F6", x"C9", x"EE", x"F2", x"F2", x"F3", x"D7", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"C5", x"EE", x"EE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"E9", x"CE", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"CE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"E9", x"EE", x"C9", x"EE", x"F2", x"F7", x"D7", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"C9", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C5", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"E9", x"F2", x"EE", x"EE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"C9", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"C5", x"E9", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"C9", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C5", x"ED", x"EE", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"C9", x"CE", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C5", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C5", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"C9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"E9", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"C9", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"EA", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"EE", x"EE", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"E9", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"CE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"E9", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EA", x"F2", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"F2", x"EA", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EA", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D2", x"F2", x"EE", x"C9", x"F2", x"EE", x"C9", x"C9", x"CD", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"E9", x"C5", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"D1", x"ED", x"D1", x"F1", x"ED", x"D1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"ED", x"F1", x"ED", x"C9", x"EE", x"F2", x"F2", x"EE", x"C9", x"D2", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"CD", x"CD", x"D1", x"F1", x"F5", x"F6", x"F1", x"F6", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"D1", x"F1", x"F1", x"C9", x"EE", x"F2", x"EE", x"EA", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"CD", x"CD", x"ED", x"F1", x"F5", x"F1", x"F1", x"F5", x"F5", x"F6", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"AC", x"CD", x"F1", x"F1", x"F1", x"CD", x"C9", x"CD", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"CD", x"ED", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"FB", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D6", x"F1", x"F1", x"F5", x"F5", x"F5", x"F1", x"CD", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"F5", x"F5", x"F1", x"F5", x"F5", x"F1", x"D1", x"FB", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"D1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"CD", x"D1", x"FB"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CC", x"F5", x"F1", x"F1", x"D1", x"F1", x"D1", x"D1", x"CD", x"D1", x"D6"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F1", x"F1", x"F1", x"F5", x"F1", x"F1", x"D1", x"F5", x"CD", x"F1", x"D1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AC", x"F5", x"F1", x"AD", x"D1", x"CD", x"F1", x"CD", x"D1", x"D2", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"CD", x"D1", x"F5", x"CD", x"F5", x"F1", x"F6", x"F5", x"F1", x"F6", x"F5", x"F1", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"F5", x"F6", x"D1", x"CC", x"CD", x"AC", x"B1", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"88", x"CD", x"CD", x"A8", x"CD", x"A8", x"CD", x"CD", x"AD", x"D1", x"F1", x"CC", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"CD", x"CD", x"CD", x"AD", x"AD", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"D6", x"DA", x"DA", x"D6", x"DA", x"D6", x"FA", x"D6", x"D6", x"DA", x"D6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B1", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF")
);
constant PinkHitted_bmp: PinkHitted_bmp_array := (
("000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000"),
("000000111111111000000011000000000000000000000000000000000000000"),
("000001111111111100000011100000000000000000000000000000000000000"),
("000011111111111110000101100000000000000000000000000000000000000"),
("000011111111111111000111100000000000000000000000000000000000000"),
("000111111111111111111111111000000000000000000000000000000000000"),
("000111111111111111111111111000000000000000000000000000000000000"),
("011111111111111111111111110000000000000000000111111110000000000"),
("011111111111111111111111110010000000000000000111111111000000000"),
("010001111111111111111111111111110000000000000011111111100000000"),
("000000111111111111111111111111110000000001111111111111110000000"),
("000000111111111111111111111111110000000001111111111111110000000"),
("000000001111111111111111111111111100000000111111111111110000000"),
("000000011111111111111111111111111100000000011111111111100000000"),
("000000011111111111111111111111111110000000011111111111100000000"),
("000001111111111111111111111111111111100001111111111111000000000"),
("000011111111111111111111111111111111110011111111111110000000000"),
("001111111111111111111111111111111111111111111111111100000000000"),
("001111111111111111111111111111111111111111111111111000000000000"),
("001111111111111111111111111111111111111111111111110000000000000"),
("001111111111111111111111111111111111111111111111000000000000000"),
("001111111111111111111111111111111111111111111110000000000000000"),
("001111111111111111111111111111111111111111111100000000000000000"),
("001111111111111111111111111111111111111111111000000000000000000"),
("000111111111111111111111111111111111111111110000000000000000000"),
("000011111111111111111111111111111111111111000000000000000000000"),
("000000111111111111111111111111111111111111100000000000000000000"),
("000000011111111111111111111111111111111111110000000000000000000"),
("000000001111111111111111111111111111111111110000000000000000000"),
("000000000111111111111111111111111111111111110000000000000000000"),
("000000000111111111111111111111111111111111110000000000000000000"),
("000000000011111111111111111111111111111111110000000000000000000"),
("000000000001111111111111111111111111111111111000000000000000000"),
("000000000000001111111111111111111111111111111100000000000000000"),
("000000000000000011111111111111111111111111111000000000000000000"),
("000000000000000011111111111111111111111111111000000000000000000"),
("000000000000000011111111111111111111111111111100000000000000000"),
("000000000000000011111111111111111111111111111110000000000000000"),
("000000000000000011111111111111111111111111111111000000000000000"),
("000000000000000011111111111111111111111111111111000000000000000"),
("000000000000000001111111111111111111111111111111100000000000000"),
("000000000000000000111111111111111111111111111111110000000000000"),
("000000000000000000111111111111111111111111111111111000000000000"),
("000000000000000000111111111111111111111111111111111000000000000"),
("000000000000000000111111111111111111111111111111111100000000000"),
("000000000000000000111111111111111111111111111111111110000000000"),
("000000000000000000111111111111111111111111111111111111000000000"),
("000000000000000000111111111111111101111111111111111111000000000"),
("000000000000000000011111111111111100111111111111111111100000000"),
("000000000000000000011111111111111100111111111111111111100000000"),
("000000000000000000011111111111111100011111111111111111100000000"),
("000000000000000001111111111111111100001111111111111111110000000"),
("000000000000000001111111111111111100000011111111111111110000000"),
("000000000000000001111111111111111100000011111111111111110000000"),
("000000000000000011111111111111111100000011111111111111110000000"),
("000000000000000011111111111111111100000011111111111111111000000"),
("000000000000000111111111111111111000000001111111111111111000000"),
("000000000000000111111111111111110000000001111111111111111000000"),
("000000000000000111111111111111110000000000111111111111111000000"),
("000000000000001111111111111111100000000000111111111111111100000"),
("000000000000001111111111111111000000000000011111111111111100000"),
("000000000000011111111111111111000000000000001111111111111110000"),
("000000000000011111111111111110000000000000000111111111111110000"),
("000000000000011111111111111100000000000000000111111111111110000"),
("000000000000111111111111111000000000000000000111111111111100000"),
("000000000000011111111111111000000000000000000011111111111000000"),
("000000000000001111111111111000000000000000000000001111111100000"),
("000000000000001111111111111000000000000000000000011111111110000"),
("000000000000001111111111000000000000000000000000011111111111000"),
("000000000000011111111110000000000000000000000000001111111111100"),
("000000000000111111111100000000000000000000000000000111111111110"),
("000000000000111111111100000000000000000000000000000111111111111"),
("000000000001111111111110000000000000000000000000000111111111111"),
("000000000001111111111111000000000000000000000000000111111111110"),
("000000000001111111111111110000000000000000000000000011111111100"),
("000000000000111111111111110000000000000000000000000001111110000"),
("000000000000111111111111100000000000000000000000000000111100000")
);
constant PinkDead_X_size : integer := 115;
constant PinkDead_Y_size : integer := 83;
type PinkDead_color_array is array(0 to PinkDead_Y_size - 1 , 0 to PinkDead_X_size - 1) of std_logic_vector(7 downto 0);
type PinkDead_bmp_array is array(0 to PinkDead_Y_size - 1 , 0 to PinkDead_X_size - 1) of std_logic;
constant PinkDead_colors: PinkDead_color_array := (
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F6", x"F6", x"F5", x"F5", x"F5", x"D1", x"F6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F6", x"F5", x"F1", x"F5", x"F5", x"F6", x"F5", x"D1", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F6", x"F7", x"FB", x"FB", x"F7", x"F7", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F6", x"FA", x"FA", x"F5", x"F6", x"F6", x"F6", x"F5", x"F6", x"F5", x"F6", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EA", x"CD", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F5", x"F6", x"F5", x"FA", x"FA", x"FA", x"F6", x"F6", x"FA", x"F6", x"F6", x"F5", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F5", x"F5", x"F1", x"D1", x"D1", x"F1", x"F6", x"FA", x"D5", x"CD", x"D1", x"D1", x"D1", x"D1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"FA", x"FA", x"FA", x"F5", x"F1", x"CD", x"CD", x"F1", x"AD", x"84", x"60", x"40", x"40", x"60", x"60", x"40", x"64", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F1", x"F5", x"F5", x"F6", x"F6", x"F5", x"F1", x"AD", x"84", x"40", x"60", x"40", x"40", x"60", x"60", x"40", x"60", x"64", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"C9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"44", x"24", x"24", x"44", x"24", x"64", x"F2", x"D6", x"F2", x"CD", x"40", x"60", x"60", x"60", x"60", x"60", x"40", x"60", x"60", x"40", x"8D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"CE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"C9", x"EE", x"EE", x"EE", x"C9", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"C9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"8E", x"CE", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"68", x"FF", x"FF", x"FB", x"F2", x"F2", x"F2", x"CE", x"FB", x"FF", x"F6", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"EE", x"C9", x"E9", x"EE", x"C9", x"C9", x"E9", x"EE", x"EE", x"EE", x"EE", x"EA", x"EE", x"EE", x"C5", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B2", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"89", x"A9", x"40", x"40", x"60", x"60", x"40", x"40", x"40", x"40", x"60", x"88", x"FB", x"F2", x"EE", x"EE", x"F2", x"EE", x"C9", x"D2", x"F6", x"C9", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"EE", x"C5", x"C9", x"C9", x"C5", x"C9", x"EE", x"C9", x"EE", x"EE", x"E9", x"EE", x"EE", x"CD", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D1", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"69", x"CD", x"84", x"60", x"40", x"40", x"60", x"60", x"60", x"60", x"60", x"84", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"C9", x"C5", x"C9", x"C9", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"EE", x"C9", x"C5", x"C5", x"C5", x"C5", x"C9", x"C9", x"C9", x"ED", x"EE", x"C9", x"E9", x"EE", x"C9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F5", x"69", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"69", x"8E", x"F2", x"F2", x"A9", x"40", x"40", x"40", x"60", x"40", x"60", x"60", x"60", x"84", x"F2", x"F2", x"D7", x"F2", x"EE", x"F2", x"D2", x"C9", x"EE", x"EE", x"C9", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"C5", x"C5", x"EE", x"C9", x"C9", x"C9", x"C9", x"EE", x"EE", x"C9", x"C9", x"EE", x"EE", x"C9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F6", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"D7", x"F2", x"F7", x"F6", x"CD", x"64", x"40", x"40", x"60", x"40", x"60", x"60", x"40", x"64", x"EE", x"EE", x"EE", x"EE", x"F2", x"D7", x"F7", x"CE", x"CE", x"C9", x"C9", x"C5", x"C9", x"C9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C5", x"C9", x"EE", x"EE", x"EE", x"EE", x"CE", x"EE", x"ED", x"E9", x"E9", x"EA", x"E9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"D1", x"F6", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"F5", x"F6", x"69", x"24", x"24", x"24", x"24", x"24", x"24", x"45", x"D2", x"D7", x"F2", x"F7", x"F7", x"F6", x"F5", x"CD", x"64", x"60", x"64", x"64", x"64", x"64", x"64", x"D1", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"EE", x"F6", x"D7", x"F2", x"E9", x"C9", x"C9", x"C9", x"C9", x"C9", x"C9", x"EE", x"ED", x"E9", x"C5", x"C9", x"ED", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"C9", x"EE", x"ED", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"FA", x"D1", x"D1", x"CD", x"CD", x"DA", x"DA", x"FA", x"F5", x"FA", x"B2", x"AD", x"F7", x"F7", x"F7", x"F2", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F5", x"D1", x"CD", x"F1", x"F6", x"F6", x"FA", x"F6", x"F6", x"F6", x"D1", x"B2", x"F2", x"F7", x"F7", x"F2", x"F7", x"F7", x"EE", x"F7", x"F7", x"F2", x"EE", x"F2", x"F2", x"EE", x"C9", x"C9", x"C9", x"C9", x"C9", x"C5", x"C5", x"C9", x"C9", x"E9", x"C9", x"E9", x"EE", x"CD", x"C9", x"C9", x"C9", x"E9", x"C5", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F6", x"D6", x"F6", x"F6", x"F6", x"D1", x"AC", x"CD", x"AD", x"F6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F3", x"F2", x"F2", x"F2", x"F7", x"D7", x"F7", x"F1", x"C9", x"CD", x"F1", x"F5", x"F1", x"F6", x"F1", x"F5", x"D1", x"88", x"20", x"65", x"CE", x"F7", x"EE", x"D7", x"F7", x"EE", x"F7", x"F7", x"F2", x"EE", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"C9", x"E9", x"C9", x"C9", x"C9", x"C9", x"C9", x"C9", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"AD", x"F5", x"AD", x"D6", x"AD", x"FA", x"D1", x"F6", x"F6", x"CD", x"CD", x"D2", x"F7", x"D7", x"F7", x"F2", x"F7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F3", x"CE", x"CD", x"F5", x"F1", x"CD", x"F5", x"D1", x"CD", x"AD", x"D2", x"AE", x"44", x"20", x"69", x"CE", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F2", x"F7", x"F7", x"D7", x"F7", x"D7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D2", x"EE", x"EE", x"D2", x"D2", x"F2", x"EE", x"EE", x"F6", x"FF", x"FF", x"FB", x"FB", x"FB", x"F7", x"F7", x"D6", x"F7", x"F6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"AC", x"D1", x"D1", x"F6", x"D1", x"F6", x"D2", x"AC", x"D1", x"F5", x"F1", x"CD", x"ED", x"F7", x"CE", x"F7", x"AD", x"44", x"AE", x"69", x"65", x"CE", x"F2", x"F2", x"EE", x"EE", x"F2", x"F7", x"EE", x"EE", x"D7", x"EE", x"CD", x"D1", x"CD", x"A8", x"CD", x"64", x"20", x"A9", x"F7", x"F7", x"CE", x"20", x"00", x"65", x"D2", x"F7", x"F7", x"F2", x"F7", x"F7", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"AC", x"D6", x"84", x"AC", x"AD", x"44", x"D1", x"F6", x"F5", x"F1", x"F6", x"F5", x"F1", x"ED", x"F2", x"F7", x"45", x"89", x"89", x"D1", x"F1", x"CD", x"F1", x"F5", x"F6", x"FA", x"F6", x"F5", x"F1", x"ED", x"D2", x"C9", x"F2", x"EE", x"EE", x"F2", x"EE", x"EE", x"A9", x"00", x"00", x"24", x"F2", x"F7", x"F2", x"40", x"00", x"00", x"69", x"F7", x"F2", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F3", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"FA", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FB", x"B1", x"FF", x"88", x"88", x"AC", x"48", x"92", x"F1", x"F5", x"FA", x"F5", x"D1", x"F5", x"F2", x"F7", x"CE", x"D2", x"24", x"69", x"FA", x"FA", x"F1", x"F1", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F1", x"CD", x"C9", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"C9", x"64", x"00", x"20", x"F2", x"F7", x"EE", x"40", x"00", x"00", x"64", x"C9", x"A9", x"C5", x"A9", x"AE", x"AE", x"AE", x"AE", x"B2", x"F6", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"FB", x"D1", x"CD", x"F1", x"F1", x"CD", x"CD", x"D1", x"F1", x"F5", x"F5", x"F1", x"CD", x"F1", x"F1", x"D2", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FB", x"B1", x"FF", x"88", x"AC", x"B1", x"00", x"AD", x"F1", x"CD", x"D1", x"CC", x"CC", x"CD", x"F2", x"B2", x"24", x"44", x"8D", x"FA", x"FA", x"FA", x"F5", x"F1", x"F6", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F5", x"F1", x"D1", x"F6", x"FA", x"FA", x"FA", x"F6", x"F1", x"CD", x"88", x"00", x"20", x"E9", x"EE", x"C9", x"44", x"40", x"40", x"40", x"40", x"60", x"60", x"40", x"40", x"60", x"40", x"40", x"64", x"F1", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"CD", x"CD", x"D1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F5", x"F6", x"D1", x"FB"),
( x"FF", x"FF", x"FF", x"FF", x"FB", x"B1", x"FF", x"88", x"AC", x"AD", x"20", x"AD", x"F5", x"88", x"AC", x"F5", x"D1", x"A8", x"F2", x"89", x"00", x"00", x"D1", x"F6", x"FA", x"FA", x"F6", x"F5", x"F5", x"F6", x"F6", x"FA", x"F6", x"F5", x"F1", x"F1", x"F5", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F5", x"F1", x"F1", x"AD", x"AD", x"F1", x"ED", x"A8", x"60", x"60", x"60", x"60", x"60", x"40", x"40", x"40", x"60", x"60", x"60", x"40", x"64", x"CD", x"D1", x"F1", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"CD", x"CD", x"ED", x"F1", x"F5", x"F5", x"F5", x"F1", x"F5", x"F5", x"F1", x"F1", x"D1", x"F1", x"CD", x"FB"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"D6", x"AD", x"88", x"88", x"88", x"AC", x"D1", x"88", x"AC", x"D5", x"A8", x"88", x"D2", x"85", x"00", x"00", x"D5", x"FA", x"FA", x"F6", x"F5", x"F5", x"F1", x"F6", x"FA", x"FA", x"F6", x"F5", x"F5", x"F6", x"F6", x"FA", x"FA", x"F6", x"FA", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"FA", x"FA", x"FA", x"88", x"40", x"60", x"60", x"40", x"40", x"40", x"40", x"60", x"60", x"40", x"40", x"40", x"64", x"F1", x"CD", x"CD", x"F2", x"F2", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F3", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F6", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F1", x"F1", x"ED", x"F1", x"F1", x"F5", x"F5", x"F1", x"F5", x"F5", x"F5", x"F1", x"F5", x"F1", x"D1", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"DB", x"DA", x"FA", x"DA", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"AD", x"EE", x"CE", x"F2", x"AD", x"20", x"00", x"D5", x"FA", x"FA", x"FA", x"F6", x"F5", x"F1", x"F5", x"F5", x"F6", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F6", x"F5", x"F6", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"88", x"60", x"40", x"60", x"60", x"40", x"40", x"60", x"60", x"60", x"60", x"60", x"40", x"64", x"F1", x"F1", x"A8", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"F1", x"CD", x"D1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F5", x"F1", x"F6", x"FF"),
( x"FF", x"FF", x"FB", x"D2", x"88", x"84", x"88", x"88", x"88", x"88", x"84", x"88", x"88", x"88", x"88", x"84", x"C9", x"F2", x"F2", x"EE", x"89", x"20", x"8D", x"F6", x"F6", x"F6", x"F5", x"D1", x"F1", x"F5", x"FA", x"FA", x"FA", x"F6", x"F5", x"F5", x"F1", x"F5", x"F6", x"F6", x"FA", x"FA", x"FA", x"FA", x"F6", x"F6", x"F6", x"F1", x"F1", x"F1", x"88", x"40", x"60", x"60", x"60", x"40", x"40", x"60", x"60", x"40", x"60", x"40", x"40", x"64", x"D1", x"CD", x"CD", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"C9", x"D1", x"D1", x"CD", x"D2", x"D1", x"CD", x"F1", x"F1", x"F1", x"F5", x"F1", x"F1", x"D1", x"CD", x"D6", x"FF"),
( x"FF", x"D6", x"88", x"84", x"88", x"A8", x"A8", x"88", x"88", x"84", x"84", x"84", x"88", x"64", x"88", x"84", x"C9", x"EE", x"EA", x"EE", x"EE", x"89", x"20", x"8D", x"F5", x"F5", x"CD", x"AD", x"CD", x"F1", x"F6", x"F6", x"F6", x"F5", x"F1", x"F1", x"F1", x"F6", x"F6", x"F6", x"F6", x"F6", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"A8", x"60", x"60", x"60", x"40", x"64", x"40", x"40", x"40", x"40", x"40", x"40", x"40", x"A9", x"D1", x"A8", x"C5", x"C9", x"E9", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"D6", x"DA", x"FF", x"FF", x"D6", x"CD", x"CD", x"F1", x"F1", x"F1", x"D1", x"F1", x"D1", x"FF", x"FF"),
( x"FF", x"AD", x"88", x"D6", x"B1", x"88", x"88", x"D6", x"D6", x"88", x"88", x"88", x"88", x"88", x"84", x"88", x"84", x"C9", x"F2", x"F2", x"EE", x"EE", x"A9", x"89", x"64", x"44", x"44", x"A9", x"CD", x"CD", x"D1", x"F1", x"F1", x"F1", x"D1", x"D1", x"F6", x"F5", x"F6", x"F5", x"F1", x"F5", x"F6", x"F6", x"F5", x"F5", x"F5", x"F1", x"CD", x"D6", x"FA", x"64", x"40", x"60", x"60", x"40", x"60", x"64", x"A8", x"A8", x"A8", x"A8", x"A8", x"F1", x"D1", x"88", x"D6", x"FB", x"FB", x"FB", x"FB", x"FB", x"EE", x"C9", x"C9", x"C9", x"E9", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"E9", x"C9", x"C9", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"CD", x"F1", x"F5", x"CD", x"CD", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"AD", x"D1", x"FF", x"FB", x"B1", x"AD", x"B1", x"D6", x"8C", x"AC", x"AC", x"AD", x"FB", x"B2", x"D6", x"FB", x"FB", x"F6", x"FF", x"FF", x"F7", x"F2", x"CE", x"CE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D6", x"D6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"D6", x"FB", x"FF", x"FF", x"FF", x"FB", x"8D", x"8D", x"8D", x"8D", x"B1", x"FB", x"FF", x"FF", x"D6", x"D6", x"F6", x"F6", x"D6", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"FB", x"FB", x"C9", x"C9", x"C9", x"C9", x"E9", x"C9", x"F2", x"FB", x"FB", x"EE", x"C9", x"EE", x"EE", x"EE", x"C9", x"EE", x"FB", x"FB", x"FB", x"FB", x"FB", x"F6", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"D1", x"D1", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
);
constant PinkDead_bmp: PinkDead_bmp_array := (
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000001111111111100000000000000000000000001111111110000000000000000000000000000000000"),
("0000000000000000000000000000000000111111111111100000000000000000000000111111111111000000000000000000000000000000000"),
("0000000000000000000000000000000001111111111111100000000000000000000011111111111111100000000000000000000000000000000"),
("0000000000000000000000000000000111111111111111110000000000000000001111111111111111110000000000000000000000000000000"),
("0000000000000000000000000000001111111111111111110000000000000001111111111111111111111100000000000000000000000000000"),
("0000000000000000000000000000011111111111111111110000000000000011111111111111111111111100000000000000000000000000000"),
("0000000000000000000000000001111111111111111111111000000000001111111111111111111111111100000000000000000000000000000"),
("0000000000000000000000000111111111111111111111111001111110111111111111111111111111111100000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000"),
("0000000000000000000000011111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000"),
("0000000000000000000000011111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000"),
("0000000000000000000000011111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000"),
("0000000000000011111000011111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000"),
("0000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000"),
("0000000000011111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000"),
("0000000001111111111111111111111111111111111111111111111111111111111111111111111111110011111111100000000000000000000"),
("0000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011110000"),
("0000110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("0000110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("0000110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("0000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("0000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("0011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111100"),
("0111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111000"),
("0011011111111111111100111110000000000111111111110001111111001111110000001111111111111111111111111111000000001110000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);
constant PinkIdle_X_size : integer := 59;
constant PinkIdle_Y_size : integer := 83;
type PinkIdle_color_array is array(0 to PinkIdle_Y_size - 1 , 0 to PinkIdle_X_size - 1) of std_logic_vector(7 downto 0);
type PinkIdle_bmp_array is array(0 to PinkIdle_Y_size - 1 , 0 to PinkIdle_X_size - 1) of std_logic;
constant PinkIdle_colors: PinkIdle_color_array := (
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"8D", x"AD", x"8D", x"AD", x"AD", x"8D", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"8D", x"68", x"64", x"64", x"64", x"64", x"64", x"64", x"88", x"8D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B2", x"64", x"64", x"64", x"64", x"88", x"68", x"64", x"68", x"88", x"64", x"68", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"88", x"64", x"64", x"64", x"64", x"64", x"68", x"68", x"64", x"88", x"64", x"64", x"8D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"64", x"64", x"64", x"64", x"64", x"CC", x"88", x"88", x"D1", x"68", x"64", x"64", x"68", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"D6", x"8D", x"64", x"68", x"64", x"64", x"64", x"A8", x"68", x"D1", x"F5", x"D1", x"64", x"88", x"68", x"8D", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"68", x"88", x"84", x"64", x"AC", x"AC", x"64", x"88", x"44", x"00", x"48", x"F1", x"F6", x"D1", x"AD", x"20", x"6D", x"8D", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"64", x"84", x"64", x"64", x"D1", x"F5", x"88", x"AC", x"D1", x"88", x"00", x"44", x"D1", x"D1", x"24", x"49", x"DF", x"89", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F7", x"FB", x"CE", x"C9", x"D2", x"D2", x"88", x"C5", x"84", x"CD", x"AD", x"D1", x"AC", x"D1", x"F5", x"D6", x"44", x"24", x"8D", x"48", x"25", x"FF", x"DB", x"8D", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"D6", x"F6", x"D6", x"D6", x"D6", x"CE", x"C9", x"D2", x"D2", x"CE", x"C5", x"A9", x"CD", x"C9", x"CD", x"D5", x"D1", x"AD", x"CD", x"F1", x"F6", x"F6", x"D5", x"D1", x"F5", x"D1", x"D1", x"FB", x"8D", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"D1", x"F1", x"D1", x"68", x"44", x"AE", x"D7", x"D2", x"D2", x"CE", x"CE", x"D2", x"CA", x"CD", x"F1", x"F6", x"F5", x"D1", x"AC", x"F1", x"F5", x"F5", x"D1", x"AD", x"AD", x"D1", x"D6", x"DB", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"F5", x"F6", x"D5", x"F5", x"69", x"00", x"89", x"D2", x"CE", x"CE", x"AE", x"D2", x"CE", x"A9", x"D1", x"F5", x"F6", x"D5", x"D1", x"AD", x"CD", x"D5", x"D1", x"AD", x"D1", x"AD", x"88", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"D5", x"F5", x"F5", x"F6", x"F6", x"D5", x"D1", x"8E", x"D2", x"CE", x"CE", x"CD", x"D2", x"CE", x"A8", x"CD", x"CD", x"D1", x"F5", x"F1", x"CD", x"AD", x"A9", x"CD", x"D1", x"D1", x"AD", x"AC", x"88", x"A9", x"C9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"F5", x"F6", x"F5", x"D6", x"F6", x"F5", x"68", x"69", x"D2", x"C9", x"C9", x"CE", x"D3", x"89", x"CD", x"AC", x"CC", x"CD", x"D1", x"CD", x"D1", x"AD", x"CD", x"AD", x"AD", x"A8", x"84", x"89", x"88", x"C9", x"D2", x"D2", x"C9", x"D7", x"CA", x"CE", x"D2", x"EE", x"EE", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F5", x"D6", x"F6", x"D5", x"F5", x"D1", x"69", x"65", x"CE", x"A9", x"CE", x"D7", x"CE", x"24", x"48", x"8D", x"AD", x"A8", x"AD", x"CD", x"D1", x"AD", x"AD", x"D1", x"F1", x"CD", x"D2", x"D6", x"D2", x"CA", x"D2", x"D2", x"D2", x"D2", x"6D", x"69", x"65", x"85", x"ED", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"CD", x"F1", x"F1", x"F1", x"F1", x"D1", x"D1", x"B1", x"CD", x"A9", x"A9", x"D2", x"D2", x"69", x"20", x"00", x"04", x"8D", x"88", x"44", x"68", x"CD", x"D1", x"D1", x"AD", x"C9", x"D2", x"D7", x"D2", x"CA", x"D2", x"D6", x"8D", x"49", x"44", x"20", x"48", x"68", x"AD", x"D1", x"A9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"CD", x"F1", x"D1", x"D1", x"D1", x"F1", x"F5", x"F6", x"D5", x"D1", x"A9", x"D2", x"CE", x"44", x"00", x"00", x"00", x"20", x"20", x"20", x"20", x"68", x"D1", x"AD", x"88", x"68", x"D6", x"D2", x"C9", x"CE", x"D2", x"D7", x"AD", x"65", x"20", x"8D", x"F6", x"D6", x"F6", x"D5", x"CD", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"F1", x"CD", x"F1", x"D5", x"F1", x"F6", x"F5", x"D6", x"F6", x"D5", x"AD", x"D2", x"65", x"00", x"00", x"00", x"20", x"40", x"20", x"20", x"20", x"20", x"68", x"D1", x"D1", x"AC", x"88", x"C9", x"CE", x"D2", x"D2", x"CE", x"AD", x"A9", x"AD", x"D5", x"D5", x"F6", x"D6", x"F5", x"F1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"F1", x"D1", x"F1", x"D5", x"F1", x"D1", x"D1", x"D1", x"F5", x"D5", x"A9", x"CD", x"44", x"20", x"20", x"40", x"40", x"40", x"20", x"40", x"40", x"20", x"49", x"D1", x"D1", x"8D", x"88", x"C9", x"C9", x"D6", x"D2", x"89", x"20", x"24", x"B1", x"D5", x"F6", x"F5", x"D5", x"F1", x"F1", x"AD", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"D1", x"F6", x"F6", x"F5", x"D5", x"D1", x"D1", x"AD", x"AC", x"AD", x"CD", x"88", x"64", x"20", x"20", x"20", x"40", x"40", x"40", x"40", x"20", x"40", x"20", x"68", x"F1", x"D1", x"AD", x"AD", x"AE", x"D2", x"D2", x"D7", x"AD", x"48", x"AD", x"D5", x"F6", x"D1", x"D1", x"D1", x"F1", x"D1", x"AD", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"D1", x"F5", x"D5", x"F6", x"D6", x"D1", x"CD", x"AD", x"AC", x"40", x"40", x"40", x"40", x"20", x"20", x"40", x"20", x"40", x"40", x"20", x"20", x"AD", x"D5", x"D1", x"AD", x"AD", x"D7", x"D2", x"D3", x"D2", x"69", x"44", x"D1", x"D1", x"F1", x"D1", x"D1", x"F1", x"F1", x"D1", x"A8", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"AD", x"AD", x"F1", x"D5", x"D6", x"F6", x"D5", x"D5", x"D1", x"F5", x"D1", x"40", x"40", x"40", x"40", x"20", x"20", x"20", x"40", x"20", x"20", x"40", x"24", x"D1", x"AD", x"AD", x"D0", x"CD", x"D2", x"CD", x"D2", x"D7", x"B2", x"45", x"88", x"CD", x"D1", x"F1", x"CD", x"CD", x"CD", x"AD", x"A8", x"AD", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"88", x"D1", x"F5", x"D5", x"F5", x"F6", x"D5", x"F5", x"D5", x"D1", x"44", x"40", x"20", x"40", x"40", x"20", x"20", x"40", x"64", x"AD", x"24", x"24", x"88", x"89", x"CD", x"CD", x"D6", x"D2", x"C9", x"CE", x"D2", x"CE", x"C9", x"89", x"88", x"A8", x"AC", x"CD", x"CD", x"CC", x"AD", x"AD", x"D1", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"8D", x"CD", x"D1", x"F1", x"F5", x"D5", x"F5", x"D5", x"D5", x"D1", x"89", x"44", x"40", x"20", x"20", x"40", x"40", x"40", x"AD", x"D2", x"CE", x"C9", x"AE", x"D6", x"D6", x"D7", x"D7", x"D2", x"C9", x"CA", x"CE", x"EE", x"A9", x"AD", x"D1", x"D1", x"CC", x"CD", x"CD", x"F1", x"D1", x"CD", x"D1", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AC", x"D1", x"CD", x"D1", x"D1", x"F1", x"D1", x"D1", x"CD", x"CD", x"CD", x"64", x"40", x"20", x"20", x"64", x"8D", x"D2", x"CE", x"CD", x"AE", x"D7", x"D7", x"D6", x"D7", x"D2", x"CE", x"CE", x"CE", x"C9", x"CE", x"A9", x"AC", x"F1", x"D1", x"D1", x"D1", x"D1", x"D1", x"D1", x"CD", x"D1", x"CD", x"89", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"F1", x"CD", x"D1", x"D1", x"F1", x"F1", x"F1", x"D1", x"D1", x"CD", x"AD", x"89", x"20", x"44", x"C9", x"D2", x"CE", x"CA", x"CD", x"D7", x"D7", x"D7", x"D7", x"D6", x"D2", x"CE", x"CE", x"CE", x"CE", x"C9", x"A5", x"88", x"CD", x"D1", x"AD", x"CD", x"CD", x"D1", x"D1", x"F1", x"D1", x"D1", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"D1", x"CD", x"D1", x"D1", x"D1", x"CD", x"AC", x"88", x"A9", x"CD", x"CD", x"C9", x"24", x"85", x"CE", x"CE", x"CE", x"C9", x"D2", x"D6", x"D6", x"D6", x"D2", x"CE", x"CE", x"CE", x"CE", x"CE", x"EE", x"AD", x"88", x"A9", x"A8", x"AD", x"AD", x"CD", x"D1", x"D1", x"D1", x"F1", x"F1", x"D5", x"D1", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"A9", x"8D", x"8D", x"8D", x"AD", x"88", x"A9", x"CD", x"A5", x"CE", x"CE", x"C9", x"A5", x"A5", x"CE", x"CE", x"C9", x"CD", x"CE", x"CE", x"CE", x"EE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CD", x"AD", x"D1", x"B1", x"B1", x"88", x"88", x"44", x"20", x"20", x"40", x"B1", x"D1", x"F1", x"D1", x"CD", x"B2", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"A9", x"C9", x"CE", x"C5", x"C9", x"CD", x"CE", x"C9", x"C9", x"C9", x"C9", x"A9", x"C9", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CD", x"B1", x"AD", x"88", x"44", x"24", x"20", x"20", x"20", x"20", x"20", x"20", x"88", x"CC", x"CD", x"AC", x"8D", x"FB", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"C9", x"CD", x"C9", x"C9", x"C9", x"C9", x"CE", x"CE", x"C9", x"A9", x"A9", x"C9", x"C9", x"CE", x"CE", x"CE", x"CE", x"CE", x"CD", x"CD", x"CE", x"CE", x"C9", x"AD", x"AD", x"D1", x"F6", x"D1", x"64", x"20", x"20", x"20", x"40", x"20", x"40", x"88", x"D1", x"CD", x"A9", x"B2", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"F7", x"C9", x"C9", x"C9", x"C9", x"C9", x"C9", x"CE", x"CE", x"CD", x"C9", x"C9", x"A9", x"A9", x"CD", x"CE", x"C9", x"CA", x"C9", x"C9", x"A9", x"D2", x"AD", x"B1", x"AD", x"D1", x"D5", x"68", x"20", x"40", x"20", x"40", x"20", x"20", x"64", x"CD", x"D1", x"AD", x"B2", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"44", x"A5", x"A9", x"A9", x"A9", x"A9", x"A9", x"CD", x"A9", x"A9", x"A9", x"A5", x"A9", x"85", x"24", x"24", x"8D", x"DB", x"DB", x"8D", x"D1", x"D1", x"D1", x"F5", x"88", x"20", x"20", x"20", x"40", x"20", x"20", x"44", x"CD", x"CC", x"88", x"B1", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"64", x"00", x"20", x"20", x"20", x"24", x"00", x"20", x"20", x"20", x"20", x"00", x"20", x"00", x"00", x"00", x"00", x"8D", x"FF", x"FF", x"D6", x"88", x"CD", x"AD", x"D1", x"D1", x"44", x"20", x"20", x"20", x"40", x"20", x"88", x"D1", x"A8", x"8D", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AE", x"C9", x"85", x"00", x"00", x"00", x"40", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"40", x"A5", x"CD", x"A9", x"DA", x"DB", x"8D", x"AD", x"B1", x"D1", x"D5", x"64", x"20", x"20", x"40", x"40", x"44", x"AD", x"88", x"8D", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"C9", x"CE", x"C9", x"85", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"44", x"44", x"44", x"A5", x"C9", x"C9", x"A9", x"C9", x"C9", x"DB", x"8D", x"68", x"AD", x"D1", x"D1", x"64", x"20", x"20", x"20", x"64", x"A8", x"B1", x"8D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"CD", x"CE", x"EE", x"C9", x"44", x"00", x"40", x"45", x"49", x"44", x"20", x"20", x"A5", x"C9", x"C9", x"C9", x"CD", x"C9", x"A9", x"A9", x"A9", x"C9", x"CE", x"DB", x"89", x"89", x"AD", x"88", x"20", x"20", x"40", x"64", x"89", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"C9", x"CE", x"CE", x"CE", x"A9", x"20", x"00", x"A9", x"CE", x"CE", x"C5", x"20", x"00", x"24", x"CD", x"CE", x"CD", x"CE", x"C9", x"A9", x"CE", x"A9", x"C9", x"D2", x"FF", x"DB", x"DF", x"FF", x"FB", x"DB", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"A5", x"C9", x"CE", x"CE", x"64", x"00", x"00", x"A9", x"C9", x"C9", x"A9", x"20", x"00", x"20", x"C9", x"CE", x"CE", x"CE", x"C9", x"A9", x"CE", x"CE", x"A9", x"A9", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"A5", x"C9", x"C9", x"C9", x"A9", x"44", x"00", x"00", x"A9", x"CE", x"C9", x"C9", x"24", x"00", x"20", x"85", x"CE", x"CE", x"CE", x"A9", x"C9", x"CD", x"A9", x"A5", x"A5", x"AE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"A5", x"CE", x"D2", x"D2", x"CA", x"A5", x"40", x"00", x"00", x"A9", x"C9", x"C9", x"CE", x"24", x"00", x"00", x"44", x"CE", x"CD", x"C9", x"C5", x"CE", x"CE", x"C9", x"C9", x"A5", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"A9", x"D2", x"D2", x"D7", x"D7", x"D2", x"C9", x"44", x"00", x"00", x"89", x"C9", x"A9", x"CE", x"24", x"00", x"00", x"44", x"A9", x"A9", x"A9", x"C9", x"CE", x"CA", x"C9", x"CE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"D2", x"D7", x"D7", x"D7", x"D7", x"D6", x"CE", x"64", x"00", x"00", x"60", x"A5", x"A5", x"A5", x"24", x"00", x"00", x"44", x"C9", x"C9", x"C9", x"CE", x"CE", x"CE", x"CE", x"C9", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"B2", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"45", x"00", x"00", x"20", x"C9", x"C9", x"CD", x"24", x"00", x"00", x"44", x"CE", x"CE", x"CE", x"CE", x"D2", x"B6", x"D2", x"CE", x"A5", x"AE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"D7", x"D7", x"D7", x"D6", x"D6", x"D7", x"D7", x"D6", x"65", x"00", x"00", x"00", x"A9", x"CE", x"CE", x"24", x"00", x"20", x"A9", x"CE", x"CE", x"D2", x"D6", x"D7", x"D7", x"D7", x"D2", x"A9", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"D6", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"69", x"00", x"00", x"40", x"A5", x"CE", x"CE", x"24", x"00", x"44", x"C9", x"CE", x"D6", x"D7", x"D6", x"D7", x"D7", x"D7", x"D7", x"D2", x"A9", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"D2", x"D7", x"D7", x"D7", x"D7", x"D7", x"D6", x"D7", x"D7", x"D3", x"45", x"20", x"65", x"A5", x"A5", x"A9", x"C9", x"69", x"20", x"A5", x"CE", x"D2", x"D7", x"D7", x"D7", x"D7", x"D7", x"B7", x"D7", x"D6", x"CE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"D2", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D6", x"D7", x"D7", x"B2", x"AD", x"CE", x"CE", x"C9", x"A5", x"A5", x"C9", x"89", x"CE", x"D2", x"D6", x"D7", x"D7", x"D6", x"D6", x"D7", x"D6", x"D7", x"D7", x"D2", x"A5", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"CE", x"CE", x"C9", x"85", x"A5", x"C9", x"C9", x"CE", x"D2", x"D7", x"D7", x"D7", x"D7", x"D7", x"D6", x"D7", x"D7", x"D7", x"D6", x"AE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"CE", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D6", x"D2", x"EE", x"C9", x"C9", x"A9", x"DB", x"CE", x"C9", x"C9", x"CE", x"D2", x"D6", x"D7", x"D7", x"D6", x"D7", x"D6", x"D7", x"D7", x"D7", x"D7", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"D2", x"D7", x"D7", x"D7", x"D6", x"D7", x"D7", x"D7", x"D7", x"D7", x"D6", x"CE", x"CE", x"A9", x"C9", x"D7", x"FF", x"D2", x"C9", x"CE", x"C9", x"D2", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"D6", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"D2", x"D2", x"CE", x"C9", x"D2", x"FF", x"FF", x"D2", x"C9", x"CE", x"C9", x"CE", x"D6", x"D7", x"D7", x"D7", x"D6", x"D7", x"D7", x"D7", x"D7", x"D7", x"CE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"D7", x"D7", x"D7", x"D7", x"D7", x"D6", x"D7", x"D2", x"CE", x"D2", x"D6", x"D2", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"A9", x"CD", x"EE", x"CE", x"D2", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D6", x"D7", x"CE", x"CE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CE", x"D6", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"C9", x"CE", x"CE", x"CE", x"D2", x"D6", x"D6", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"CE", x"D2", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CE", x"D6", x"D2", x"D2", x"D7", x"D7", x"D7", x"D7", x"D7", x"D7", x"D2", x"CE", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"A9", x"CA", x"D2", x"D7", x"D2", x"D2", x"D2", x"D6", x"D6", x"D7", x"D7", x"D7", x"D7", x"D2", x"CE", x"D6", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EE", x"D2", x"CE", x"CE", x"F2", x"D7", x"D7", x"D7", x"D2", x"D2", x"C9", x"C5", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"D2", x"D6", x"D7", x"D6", x"D2", x"D7", x"D2", x"D2", x"D2", x"D7", x"D7", x"D7", x"CE", x"D2", x"CE", x"A9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"EE", x"EE", x"EE", x"CE", x"D6", x"D7", x"D7", x"D2", x"EE", x"C9", x"AD", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"A9", x"CE", x"D2", x"D6", x"D7", x"D7", x"D7", x"D2", x"CE", x"CA", x"D2", x"D2", x"D2", x"CE", x"EE", x"CE", x"CE", x"CE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"D6", x"D2", x"EE", x"CE", x"D2", x"CD", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"EE", x"D2", x"D6", x"D7", x"D7", x"D7", x"D2", x"CE", x"C9", x"C9", x"CE", x"CE", x"EE", x"EE", x"EE", x"CE", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"C9", x"EE", x"CE", x"EE", x"EE", x"EE", x"CE", x"D2", x"D6", x"D2", x"CE", x"C9", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"CE", x"CE", x"F2", x"D6", x"D6", x"D6", x"D2", x"CE", x"CE", x"CE", x"EE", x"CE", x"CE", x"EE", x"CE", x"CE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"CE", x"EE", x"EE", x"CE", x"EE", x"EE", x"CE", x"D2", x"D2", x"CE", x"C9", x"C9", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"A9", x"CE", x"CE", x"CE", x"CE", x"EE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"CE", x"EE", x"CE", x"CE", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"CE", x"CE", x"EE", x"EE", x"EE", x"CE", x"EE", x"EE", x"EE", x"C9", x"CD", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"A5", x"C9", x"CE", x"CE", x"EE", x"CE", x"CE", x"EE", x"CE", x"EE", x"EE", x"CE", x"EE", x"CE", x"EE", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"CE", x"EE", x"CE", x"CD", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D2", x"C9", x"CE", x"CE", x"EE", x"CE", x"EE", x"EE", x"CE", x"CE", x"EE", x"EE", x"CE", x"CE", x"C9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"EE", x"EE", x"CE", x"C5", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"A5", x"C9", x"EE", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"CD", x"CE", x"CE", x"CE", x"CE", x"CE", x"EE", x"EE", x"CE", x"EE", x"EE", x"EE", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"A9", x"EE", x"CE", x"CE", x"CE", x"F2", x"EE", x"CE", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"D2", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CD", x"D2", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"CE", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"A9", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CD", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"EE", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"C9", x"A5", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C5", x"CE", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"A9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"F2", x"EE", x"EE", x"CE", x"CD", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C5", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CD", x"CD", x"AD", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CE", x"CD", x"EE", x"F2", x"CE", x"EE", x"EE", x"CE", x"EE", x"CE", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"CD", x"C9", x"CE", x"F2", x"F2", x"EE", x"EE", x"EE", x"CE", x"C9", x"AD", x"CD", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"A9", x"CD", x"C9", x"C9", x"EE", x"CD", x"CD", x"FA", x"CE", x"D7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"CA", x"D2", x"CA", x"C9", x"EE", x"CE", x"CD", x"CD", x"F1", x"D1", x"D1", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F1", x"F1", x"D1", x"ED", x"F1", x"F1", x"AD", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"A9", x"CD", x"ED", x"F1", x"F1", x"F1", x"F5", x"D1", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F1", x"F1", x"F5", x"F5", x"F1", x"F1", x"D1", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"F1", x"F1", x"F5", x"F1", x"F5", x"F1", x"F1", x"CD", x"D2", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F1", x"F5", x"F5", x"F5", x"F1", x"F5", x"F1", x"F1", x"D1", x"8C", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F5", x"D1", x"F5", x"F1", x"F5", x"F1", x"F1", x"F1", x"CD", x"D2", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F1", x"F1", x"F1", x"F5", x"F1", x"F1", x"F5", x"F1", x"D1", x"D1", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AD", x"F1", x"F1", x"F1", x"F1", x"F1", x"ED", x"F1", x"D1", x"F1", x"CD", x"CC", x"D6", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"D6", x"D6", x"D1", x"F1", x"D1", x"F1", x"F1", x"D1", x"ED", x"F1", x"F1", x"F5", x"F1", x"CD", x"A9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"F1", x"F6", x"F1", x"F1", x"CD", x"F5", x"D1", x"F1", x"D1", x"D1", x"CD", x"F1", x"AD", x"FF", x"FF"),
( x"FF", x"FF", x"D6", x"F2", x"CD", x"D1", x"D1", x"D1", x"D1", x"CD", x"F1", x"D5", x"F5", x"F1", x"F1", x"F5", x"CD", x"D6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"F1", x"F5", x"F5", x"D1", x"CD", x"D5", x"CD", x"D1", x"D1", x"88", x"AD", x"AC", x"A8", x"FB", x"FF"),
( x"FF", x"FF", x"D1", x"CD", x"CC", x"AC", x"AC", x"D1", x"F1", x"A8", x"F1", x"F5", x"F5", x"F1", x"CD", x"CD", x"8C", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"88", x"AD", x"AD", x"A8", x"D6", x"AD", x"AD", x"A8", x"AD", x"AC", x"DA", x"FF", x"FB", x"FB", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"D2", x"AD", x"AD", x"AD", x"AD", x"D1", x"D6", x"AD", x"B1", x"D1", x"CD", x"AD", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
);
constant PinkIdle_bmp: PinkIdle_bmp_array := (
("00000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000111111110000000000000000000000"),
("00000000000000000000000000001111111111000000000000000000000"),
("00000000000000000000000000011111111111100000000000000000000"),
("00000000000000000000000000011111111111110000000000000000000"),
("00000000000000000000000000111111111111111000000000000000000"),
("00000000000000000000000011111111111111111100000000000000000"),
("00000000000000000000000011111111111111111110000000000000000"),
("00000000000000000000000011111111111111111110000000000000000"),
("00000000000000000111111111111111111111101110000000000000000"),
("00000000000111111111111111111111111111111100000000000000000"),
("00000000001111111111111111111111111111111000000000000000000"),
("00000000011111111111111111111111111111000000000000000000000"),
("00000000111111111111111111111111111111111000000000000000000"),
("00000000111111111111111111111111111111111111111111000000000"),
("00000000111111111111111111111111111111111111111111000000000"),
("00000001111111111111111111111111111111111111111110000000000"),
("00000001111111111111111111111111111111111111111111000000000"),
("00000011111111111111111111111111111111111111111111100000000"),
("00000011111111111111111111111111111111111111111111100000000"),
("00000011111111111111111111111111111111111111111111100000000"),
("00000011111111111111111111111111111111111111111111100000000"),
("00000011111111111111111111111111111111111111111111110000000"),
("00000001111111111111111111111111111111111111111111111000000"),
("00000000111111111111111111111111111111111111111111111000000"),
("00000000111111111111111111111111111111111111111111111000000"),
("00000000011111111111111111111111111111111111111111111000000"),
("00000000011111111111111111111111111111111111111111111100000"),
("00000000011111111111111111111111111111111111111111111110000"),
("00000000000000111111111111111111111111111111111111111111000"),
("00000000000000011111111111111111111111111111111111111111000"),
("00000000000000001111111111111111111111111111111111111111000"),
("00000000000000000011111111111111111111111111111111111111000"),
("00000000000000000011111111111111111110011111111111111110000"),
("00000000000000000111111111111111111111111111111111111100000"),
("00000000000000001111111111111111111111111111111111111000000"),
("00000000000000001111111111111111111111111111111111110000000"),
("00000000000000011111111111111111111111110110111100000000000"),
("00000000000000011111111111111111111111111000000000000000000"),
("00000000000000111111111111111111111111111000000000000000000"),
("00000000000001111111111111111111111111111000000000000000000"),
("00000000000001111111111111111111111111110000000000000000000"),
("00000000000011111111111111111111111111111000000000000000000"),
("00000000000111111111111111111111111111111000000000000000000"),
("00000000001111111111111111111111111111111000000000000000000"),
("00000000001111111111111111111111111111111100000000000000000"),
("00000000011111111111111111111111111111111110000000000000000"),
("00000000011111111111111111111111111111111110000000000000000"),
("00000000111111111111111111111111111111111110000000000000000"),
("00000000111111111111111111111111111111111110000000000000000"),
("00000000111111111111111110111111111111111110000000000000000"),
("00000000111111111111111100111111111111111110000000000000000"),
("00000000111111111111111000011111111111111111000000000000000"),
("00000001111111111111110000011111111111111111100000000000000"),
("00000001111111111111100000001111111111111111110000000000000"),
("00000001111111111111100000001111111111111111111000000000000"),
("00000001111111111111100000000111111111111111111100000000000"),
("00000001111111111111100000000111111111111111111100000000000"),
("00000011111111111111100000000011111111111111111110000000000"),
("00000011111111111111100000000001111111111111111110000000000"),
("00000011111111111111100000000000111111111111111110000000000"),
("00000011111111111111110000000000011111111111111111000000000"),
("00000001111111111111110000000000001111111111111111000000000"),
("00000001111111111111110000000000000111111111111111100000000"),
("00000001111111111111110000000000000111111111111111111000000"),
("00000001111111111111110000000000000011111111111111111000000"),
("00000000111111111111110000000000000001111111111111110000000"),
("00000001111111111111111000000000000000111111111111110000000"),
("00000001111111111111111000000000000000111111111111111000000"),
("00000000111111111111100000000000000000011111111111111000000"),
("00000000011111111111000000000000000000001111111111111000000"),
("00000000011111111110000000000000000000000000111111111100000"),
("00000000111111111110000000000000000000000000011111111110000"),
("00000001111111111110000000000000000000000000111111111111000"),
("00000011111111111110000000000000000000000001111111111111100"),
("00001111111111111110000000000000000000000001111111111111100"),
("00111111111111111110000000000000000000000001111111111111110"),
("00111111111111111100000000000000000000000001111111111101100"),
("00011111111111110000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000")
);
constant PinkWon_X_size : integer := 66;
constant PinkWon_Y_size : integer := 83;
type PinkWon_color_array is array(0 to PinkWon_Y_size - 1 , 0 to PinkWon_X_size - 1) of std_logic_vector(7 downto 0);
type PinkWon_bmp_array is array(0 to PinkWon_Y_size - 1 , 0 to PinkWon_X_size - 1) of std_logic;
constant PinkWon_colors: PinkWon_color_array := (
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D6", x"88", x"88", x"88", x"88", x"88", x"88", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"88", x"84", x"88", x"88", x"88", x"88", x"88", x"88", x"88", x"AC", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"88", x"88", x"AC", x"88", x"88", x"88", x"88", x"AC", x"88", x"88", x"84", x"88", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"88", x"88", x"D1", x"88", x"88", x"AC", x"D1", x"A8", x"88", x"88", x"88", x"84", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"88", x"AD", x"D1", x"CD", x"AC", x"F6", x"B1", x"AD", x"88", x"CD", x"AC", x"84", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"44", x"00", x"20", x"68", x"FA", x"D6", x"24", x"44", x"44", x"20", x"88", x"88", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"44", x"64", x"88", x"44", x"F6", x"D1", x"89", x"AC", x"A8", x"68", x"B1", x"AD", x"CE", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"64", x"CC", x"AC", x"88", x"D5", x"D1", x"CD", x"D1", x"D1", x"AC", x"F5", x"D1", x"C9", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"AD", x"AD", x"D1", x"88", x"CD", x"88", x"AC", x"F5", x"FA", x"FA", x"F5", x"CD", x"CD", x"A8", x"88", x"88", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"FB", x"FB", x"AD", x"D6", x"D1", x"F1", x"A8", x"D1", x"A8", x"AD", x"CD", x"F6", x"FA", x"F5", x"F1", x"F5", x"F5", x"88", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F6", x"F2", x"EE", x"F2", x"D2", x"CD", x"A8", x"D1", x"AC", x"CD", x"CC", x"D1", x"F5", x"F1", x"CD", x"F2", x"F2", x"A8", x"88", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"EE", x"F2", x"F2", x"C5", x"84", x"64", x"88", x"AC", x"B1", x"D1", x"A8", x"F1", x"CC", x"ED", x"F6", x"F2", x"CE", x"CD", x"88", x"DA", x"FF", x"FF", x"FF", x"F6", x"F6", x"F7", x"F7", x"F2", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F2", x"F2", x"F2", x"EE", x"F7", x"CE", x"40", x"40", x"40", x"40", x"40", x"64", x"CD", x"64", x"CD", x"AD", x"8D", x"F2", x"EE", x"EE", x"EE", x"CE", x"CE", x"EE", x"EE", x"F2", x"D2", x"F2", x"F2", x"EE", x"C9", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F3", x"F7", x"F2", x"EE", x"EE", x"89", x"20", x"40", x"60", x"60", x"40", x"40", x"40", x"40", x"AD", x"24", x"65", x"F2", x"F6", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F7", x"F2", x"D2", x"C9", x"C9", x"EA", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"69", x"64", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"D2", x"F6", x"F2", x"F2", x"EE", x"D2", x"00", x"20", x"40", x"60", x"60", x"40", x"40", x"40", x"20", x"00", x"00", x"89", x"F7", x"EE", x"F7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F2", x"C9", x"40", x"44", x"C9", x"EA", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"8D", x"40", x"40", x"64", x"F5", x"F6", x"F6", x"F6", x"F6", x"F5", x"F1", x"FB", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"ED", x"EE", x"F2", x"F7", x"F2", x"D2", x"00", x"20", x"40", x"40", x"60", x"40", x"64", x"88", x"40", x"00", x"44", x"F2", x"F7", x"CE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"92", x"69", x"D5", x"F1", x"CD", x"ED", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"8D", x"40", x"40", x"40", x"40", x"64", x"F1", x"CC", x"AC", x"A8", x"A8", x"A8", x"AD", x"FB", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"EE", x"F2", x"F7", x"F2", x"D2", x"00", x"40", x"40", x"40", x"40", x"40", x"88", x"D1", x"84", x"20", x"A9", x"F2", x"F7", x"CE", x"F7", x"F7", x"F7", x"F7", x"D7", x"F2", x"F2", x"EE", x"F6", x"FA", x"FA", x"FA", x"F5", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"B6", x"40", x"64", x"AD", x"8C", x"40", x"40", x"AC", x"84", x"AD", x"D2", x"B2", x"D1", x"DB", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B2", x"AC", x"ED", x"C9", x"F2", x"F7", x"EE", x"D2", x"20", x"40", x"40", x"40", x"40", x"40", x"40", x"44", x"20", x"A9", x"F2", x"F7", x"F7", x"C9", x"F7", x"F3", x"F2", x"F7", x"F7", x"CD", x"44", x"8D", x"F6", x"FA", x"FA", x"FA", x"F6", x"F5", x"CD", x"FF", x"FF", x"FF", x"FF", x"44", x"40", x"D1", x"FA", x"F6", x"D1", x"A8", x"A8", x"A8", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"88", x"AC", x"C9", x"F2", x"F7", x"EE", x"D2", x"20", x"40", x"60", x"60", x"40", x"40", x"20", x"00", x"20", x"EE", x"F2", x"F7", x"F7", x"CE", x"F7", x"F7", x"EE", x"D2", x"CE", x"64", x"D1", x"F6", x"FA", x"FA", x"F1", x"F5", x"F5", x"F1", x"CD", x"FF", x"FF", x"FF", x"89", x"40", x"60", x"D1", x"F5", x"F1", x"F5", x"F1", x"CD", x"AD", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"F1", x"CD", x"EE", x"F7", x"EE", x"D2", x"60", x"40", x"60", x"40", x"40", x"40", x"20", x"24", x"AE", x"F7", x"F7", x"D7", x"F7", x"EE", x"F2", x"F7", x"F2", x"D2", x"A9", x"C9", x"F5", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F1", x"D6", x"FF", x"8D", x"40", x"60", x"40", x"60", x"64", x"64", x"84", x"CD", x"AC", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"CD", x"EE", x"F2", x"CD", x"CD", x"CD", x"60", x"40", x"40", x"40", x"20", x"00", x"89", x"F7", x"D7", x"EE", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"C9", x"64", x"AD", x"F1", x"F5", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F1", x"CD", x"64", x"40", x"60", x"60", x"60", x"40", x"40", x"40", x"AD", x"B2", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"CD", x"C9", x"CD", x"CD", x"F1", x"F5", x"CD", x"A8", x"88", x"64", x"40", x"44", x"D2", x"F7", x"F7", x"D2", x"F2", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"C9", x"CD", x"CD", x"F1", x"F5", x"F6", x"F5", x"FA", x"F6", x"F1", x"D1", x"CC", x"40", x"40", x"60", x"60", x"40", x"40", x"40", x"8D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F1", x"F1", x"A8", x"88", x"CD", x"F1", x"F5", x"F5", x"F5", x"F1", x"F1", x"AC", x"44", x"89", x"F7", x"D7", x"F7", x"F2", x"F2", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"A9", x"CD", x"CD", x"F1", x"F1", x"F5", x"F5", x"F6", x"F5", x"F1", x"F1", x"AD", x"40", x"40", x"60", x"60", x"40", x"40", x"40", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"CD", x"AC", x"A8", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"CD", x"64", x"64", x"D2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"C9", x"C9", x"CD", x"F1", x"F5", x"F1", x"F1", x"F1", x"F1", x"F5", x"D1", x"CD", x"CD", x"CD", x"84", x"40", x"40", x"20", x"40", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"CD", x"CC", x"A8", x"F1", x"F5", x"F5", x"F5", x"F1", x"F1", x"AD", x"84", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"CD", x"A8", x"CD", x"F1", x"F5", x"F1", x"D1", x"CD", x"CD", x"CD", x"CD", x"F1", x"F5", x"F5", x"F1", x"84", x"60", x"89", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"ED", x"CD", x"A8", x"F1", x"F1", x"F5", x"F5", x"F1", x"F1", x"A8", x"A9", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"CD", x"A8", x"CC", x"F1", x"F1", x"CD", x"CD", x"CD", x"F1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"D1", x"CC", x"A8", x"F1", x"F1", x"F1", x"F1", x"F1", x"D1", x"A8", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"AD", x"D1", x"F1", x"CD", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"CD", x"88", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"A8", x"A8", x"F1", x"ED", x"CD", x"D1", x"F1", x"CD", x"ED", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"CD", x"AD", x"AD", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"A8", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"A8", x"84", x"A8", x"C9", x"AD", x"CD", x"F2", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"C9", x"F7", x"FF", x"CD", x"CD", x"F5", x"F5", x"F1", x"F5", x"F5", x"F1", x"AC", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"E9", x"C9", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"C9", x"F2", x"FF", x"FF", x"FF", x"D1", x"F1", x"F1", x"F5", x"F5", x"F1", x"AC", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"EA", x"EE", x"C9", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"D1", x"F1", x"CD", x"AC", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"C9", x"C5", x"E9", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"C9", x"C9", x"85", x"64", x"A5", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"A8", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D7", x"44", x"20", x"40", x"44", x"A5", x"C9", x"C9", x"EE", x"CE", x"CE", x"CA", x"C9", x"C5", x"44", x"40", x"40", x"00", x"00", x"20", x"69", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"85", x"00", x"00", x"00", x"20", x"40", x"20", x"20", x"20", x"20", x"20", x"20", x"20", x"00", x"00", x"20", x"20", x"89", x"CE", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"A9", x"20", x"00", x"00", x"81", x"44", x"00", x"00", x"00", x"00", x"00", x"20", x"44", x"65", x"C9", x"EE", x"EE", x"EE", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"F2", x"F2", x"EE", x"65", x"00", x"00", x"64", x"65", x"20", x"00", x"00", x"64", x"69", x"A9", x"EE", x"F2", x"F2", x"EE", x"C9", x"E9", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"A9", x"20", x"00", x"20", x"EE", x"EE", x"A9", x"20", x"00", x"89", x"F2", x"F2", x"F2", x"EE", x"F2", x"E9", x"EE", x"E9", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F2", x"EE", x"65", x"00", x"00", x"A9", x"F2", x"EE", x"EE", x"44", x"00", x"44", x"EE", x"F2", x"F2", x"F2", x"EE", x"E9", x"EE", x"EE", x"C9", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"A9", x"00", x"00", x"00", x"EE", x"EE", x"C9", x"EE", x"44", x"00", x"40", x"CE", x"F2", x"F2", x"F2", x"EE", x"C9", x"EE", x"F2", x"C9", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"E9", x"EE", x"85", x"00", x"00", x"40", x"EE", x"EE", x"C9", x"EE", x"A5", x"20", x"00", x"89", x"F2", x"F2", x"F2", x"EE", x"EA", x"F2", x"EE", x"E9", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"EA", x"85", x"00", x"00", x"A9", x"EE", x"EE", x"EE", x"F2", x"CE", x"20", x"00", x"69", x"F2", x"EE", x"EE", x"CD", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F7", x"F2", x"A9", x"00", x"00", x"A9", x"C9", x"EE", x"EE", x"EE", x"C9", x"20", x"00", x"65", x"EE", x"EE", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"D2", x"F7", x"F2", x"85", x"00", x"00", x"A9", x"EE", x"EE", x"EE", x"EE", x"CE", x"00", x"00", x"64", x"EE", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"F7", x"F7", x"CE", x"20", x"00", x"00", x"AE", x"F2", x"EE", x"EE", x"EE", x"EE", x"20", x"00", x"65", x"EE", x"F2", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"D7", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"F7", x"F7", x"CE", x"00", x"00", x"00", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"00", x"00", x"65", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F7", x"F7", x"D7", x"69", x"00", x"00", x"44", x"CE", x"EE", x"EE", x"EE", x"C9", x"C9", x"20", x"00", x"69", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"F7", x"F7", x"D7", x"20", x"20", x"89", x"D2", x"F6", x"F2", x"EE", x"C9", x"C9", x"C5", x"65", x"00", x"69", x"F2", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F7", x"F7", x"F7", x"B2", x"B2", x"F7", x"F7", x"F7", x"F2", x"EE", x"ED", x"C9", x"C5", x"A5", x"00", x"89", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"EE", x"E9", x"C5", x"C9", x"EE", x"F3", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"EE", x"E9", x"A5", x"C9", x"EE", x"F6", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"C9", x"FB", x"E9", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"C9", x"F7", x"FF", x"C9", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"CE", x"C5", x"FF", x"FF", x"F6", x"EE", x"F7", x"D7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"E9", x"CD", x"FF", x"FF", x"FB", x"C9", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"C9", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"F7", x"F7", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EA", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"CE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"EE", x"EA", x"EE", x"C9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"EA", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"C9", x"C9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"EE", x"EE", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"C9", x"C9", x"EE", x"EE", x"EE", x"ED", x"EE", x"EE", x"EE", x"EE", x"E9", x"C5", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"C9", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F7", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"E9", x"E9", x"E9", x"EE", x"EE", x"EA", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"C9", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F7", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"EE", x"EE", x"ED", x"EE", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"C9", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C5", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"EE", x"CE", x"EE", x"EE", x"EE", x"CE", x"EE", x"EE", x"EE", x"EA", x"EE", x"E9", x"C5", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"E9", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"EE", x"CE", x"EE", x"EE", x"EA", x"EA", x"EE", x"EE", x"E9", x"EE", x"EE", x"E9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"EE", x"EE", x"ED", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"ED", x"C5", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C9", x"EE", x"EE", x"ED", x"EE", x"EA", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"C9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"EE", x"C9", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"C9", x"EE", x"EE", x"EE", x"EE", x"CE", x"EE", x"EA", x"EE", x"EA", x"EE", x"ED", x"C9", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EA", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"E9", x"EE", x"EE", x"E9", x"ED", x"EE", x"EE", x"EE", x"EE", x"EA", x"EE", x"EA", x"C5", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C5", x"C9", x"EE", x"EA", x"CE", x"EE", x"EE", x"EE", x"CD", x"ED", x"ED", x"CE", x"C9", x"C5", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"C9", x"C9", x"EE", x"E9", x"C9", x"C9", x"C9", x"CE", x"E9", x"C9", x"C9", x"C9", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"C9", x"C9", x"C9", x"C9", x"C9", x"E9", x"C9", x"C9", x"EE", x"D2", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"CE", x"EE", x"EE", x"E9", x"ED", x"F2", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"F1", x"F1", x"F1", x"ED", x"CD", x"D2", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F6", x"FF", x"F7", x"CE", x"CD", x"CD", x"ED", x"F1", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"F1", x"F1", x"D1", x"F1", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"F1", x"F1", x"ED", x"D1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"CD", x"F1", x"F1", x"F1", x"F1", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F1", x"F1", x"F1", x"ED", x"ED", x"CD", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"D1", x"F1", x"F5", x"F5", x"F1", x"F1", x"D1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"F1", x"D1", x"CD", x"CD", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"ED", x"CD", x"CD", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"CD", x"F1", x"F1", x"F5", x"F5", x"F5", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"A8", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"F5", x"F5", x"F1", x"F5", x"F5", x"F1", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F5", x"F1", x"F5", x"F1", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"F1", x"CD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"ED", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F5", x"F5", x"F5", x"F1", x"CD", x"F1", x"ED", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"CD", x"F1", x"F5", x"F5", x"F1", x"F5", x"F5", x"F5", x"F1", x"F5", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FB", x"FA", x"D1", x"AD", x"CD", x"D1", x"CD", x"F1", x"F1", x"F1", x"F5", x"F1", x"F5", x"CD", x"88", x"A8", x"A8", x"AC", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"AD", x"F1", x"F1", x"F1", x"ED", x"F1", x"F1", x"F1", x"F1", x"F1", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"CD", x"CD", x"D1", x"CD", x"F5", x"F1", x"D1", x"F6", x"F6", x"F5", x"F1", x"D1", x"CD", x"B1", x"B1", x"D6", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"F1", x"F1", x"F1", x"F5", x"D1", x"CD", x"F1", x"D1", x"D1", x"CD", x"F1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"D6", x"AD", x"AD", x"AD", x"AD", x"D1", x"AD", x"D1", x"D1", x"D1", x"D1", x"FB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"F1", x"F5", x"F6", x"F5", x"CD", x"F6", x"AD", x"D1", x"A8", x"CD", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AC", x"AD", x"AD", x"AD", x"A8", x"D6", x"CD", x"88", x"A8", x"88", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
);
constant PinkWon_bmp: PinkWon_bmp_array := (
("000000000000000000011111111110000000000000000000000000000000000000"),
("000000000000000000111111111111000000000000000000000000000000000000"),
("000000000000000001111111111111000000000000000000000000000000000000"),
("000000000000000001111111111111000000000000000000000000000000000000"),
("000000000000000001111111111111000000000000000000000000000000000000"),
("000000000000000001111111111111000000000000000000000000000000000000"),
("000000000000000001111111111111110000000000000000000000000000000000"),
("000000000000000001111111111111111000000000000000000000000000000000"),
("000000000000000011111111111111111000000000000000000000000000000000"),
("000000000000011111111111111111111100000000000000000000000000000000"),
("000000000000111111111111111111111100000000010000000000000000000000"),
("000000000000111111111111111111111110001111110000000000000000000000"),
("000000000001111111111111111111111111111111110000000000000000000000"),
("000000000001111111111111111111111111111111110000000000111100000000"),
("000000000011111111111111111111111111111111110000000011111111111110"),
("000000000111111111111111111111111111111111111000000111111111111110"),
("000000000111111111111111111111111111111111111100001111111111111100"),
("000000000111111111111111111111111111111111111100001111111111000000"),
("000000000111111111111111111111111111111111111100011111111111000000"),
("000000000111111111111111111111111111111111111110111111111110000000"),
("000000000111111111111111111111111111111111111111111111111100000000"),
("000000000111111111111111111111111111111111111111111111100000000000"),
("000000000111111111111111111111111111111111111111111111100000000000"),
("000000000111111111111111111111111111111111111111111111000000000000"),
("000000000111111111111111111111111111111111111111111110000000000000"),
("000000000011111111111111111111111111111111111111111110000000000000"),
("000000000011111111111111111111111111111111111111111100000000000000"),
("000000000011111111111111111111111111111111111111111100000000000000"),
("000000000000011111111111111111111111111101111111111000000000000000"),
("000000000000001111111111111111111111111000111111110000000000000000"),
("000000000000000111111111111111111111110000011111100000000000000000"),
("000000000000000111111111111111111111100000001110000000000000000000"),
("000000000000000011111111111111111111100000000100000000000000000000"),
("000000000000000011111111111111111111100000000000000000000000000000"),
("000000000000000111111111111111111111110000000000000000000000000000"),
("000000000000001111111111111111111111110000000000000000000000000000"),
("000000000000001111111111111111111111111000000000000000000000000000"),
("000000000000001111111111111111111111111000000000000000000000000000"),
("000000000000001111111111111111111111111000000000000000000000000000"),
("000000000000001111111111111111111111111000000000000000000000000000"),
("000000000000001111111111111111111111111000000000000000000000000000"),
("000000000000001111111111111111111111111100000000000000000000000000"),
("000000000000011111111111111111111111111100000000000000000000000000"),
("000000000000011111111111111111111111111100000000000000000000000000"),
("000000000000111111111111111111111111111100000000000000000000000000"),
("000000000000111111111111111111111111111110000000000000000000000000"),
("000000000000111111111111111111111111111110000000000000000000000000"),
("000000000000111111111111111111111111111110000000000000000000000000"),
("000000000000111111111111111111111111111110000000000000000000000000"),
("000000000000111111111111111111111111111110000000000000000000000000"),
("000000000000111111111111111111111111111111000000000000000000000000"),
("000000000000111111111111111011111111111111000000000000000000000000"),
("000000000000111111111111110011111111111111000000000000000000000000"),
("000000000000111111111111110011111111111111000000000000000000000000"),
("000000000000111111111111100001111111111111000000000000000000000000"),
("000000000000111111111111100001111111111111100000000000000000000000"),
("000000000001111111111111100000111111111111110000000000000000000000"),
("000000000001111111111111100000111111111111110000000000000000000000"),
("000000000011111111111111100000111111111111111000000000000000000000"),
("000000000111111111111111100000011111111111111000000000000000000000"),
("000000000111111111111111100000011111111111111100000000000000000000"),
("000000000111111111111111000000001111111111111100000000000000000000"),
("000000000111111111111111000000001111111111111100000000000000000000"),
("000000000111111111111111000000001111111111111100000000000000000000"),
("000000000111111111111111000000000111111111111110000000000000000000"),
("000000000111111111111110000000000111111111111110000000000000000000"),
("000000001111111111111110000000000111111111111110000000000000000000"),
("000000001111111111111110000000000011111111111110000000000000000000"),
("000000011111111111111110000000000011111111111111000000000000000000"),
("000000011111111111111110000000000011111111111110000000000000000000"),
("000000000111111111111110000000000001111111111000000000000000000000"),
("000000000001111111111000000000000001101111111000000000000000000000"),
("000000000000111111100000000000000000000111111100000000000000000000"),
("000000000001111111100000000000000000000111111110000000000000000000"),
("000000000011111111100000000000000000000111111111000000000000000000"),
("000000000111111111111000000000000000000111111111000000000000000000"),
("000000001111111111111000000000000000000111111111100000000000000000"),
("000000011111111111111000000000000000000111111111110000000000000000"),
("000001111111111111111000000000000000000111111111111000000000000000"),
("001111111111111111111000000000000000000111111111111100000000000000"),
("001111111111111111100000000000000000000111111111111110000000000000"),
("001111111111111000000000000000000000000011111111111110000000000000"),
("000000000000000000000000000000000000000001111111111100000000000000")
);
constant PinkPunch_X_size : integer := 73;
constant PinkPunch_Y_size : integer := 83;
type PinkPunch_color_array is array(0 to PinkPunch_Y_size - 1 , 0 to PinkPunch_X_size - 1) of std_logic_vector(7 downto 0);
type PinkPunch_bmp_array is array(0 to PinkPunch_Y_size - 1 , 0 to PinkPunch_X_size - 1) of std_logic;
constant PinkPunch_colors: PinkPunch_color_array := (
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"DB", x"DB", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D6", x"D6", x"D6", x"D6", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"B2", x"64", x"40", x"40", x"40", x"89", x"B6", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AD", x"84", x"84", x"84", x"84", x"84", x"64", x"8D", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"8D", x"20", x"40", x"40", x"60", x"60", x"40", x"40", x"B2", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"84", x"88", x"88", x"88", x"A8", x"84", x"88", x"88", x"88", x"88", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F1", x"D5", x"64", x"40", x"60", x"60", x"60", x"60", x"60", x"60", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"A8", x"84", x"68", x"88", x"84", x"88", x"88", x"88", x"88", x"88", x"A8", x"88", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F5", x"AD", x"20", x"40", x"40", x"40", x"60", x"40", x"40", x"60", x"89", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"64", x"88", x"88", x"88", x"88", x"CD", x"A8", x"AC", x"D1", x"A8", x"88", x"84", x"88", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"AD", x"CD", x"60", x"40", x"40", x"40", x"40", x"40", x"64", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"88", x"88", x"88", x"88", x"88", x"CD", x"8D", x"B1", x"FA", x"F6", x"CD", x"88", x"A8", x"B1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"FA", x"FA", x"F5", x"44", x"40", x"40", x"40", x"40", x"40", x"40", x"D6", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"84", x"AC", x"CC", x"88", x"A8", x"64", x"00", x"20", x"AD", x"F5", x"F6", x"CD", x"F6", x"DA", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"F5", x"AD", x"40", x"60", x"60", x"40", x"60", x"40", x"40", x"69", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AD", x"AD", x"B1", x"AD", x"AD", x"A4", x"A8", x"D5", x"F6", x"AC", x"D1", x"B1", x"24", x"68", x"00", x"89", x"F6", x"F5", x"D2", x"FF", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"64", x"40", x"60", x"60", x"60", x"40", x"40", x"40", x"89", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"89", x"A8", x"A8", x"A8", x"88", x"88", x"88", x"A8", x"A8", x"CD", x"F6", x"F1", x"F5", x"FA", x"D1", x"D6", x"44", x"24", x"AD", x"F6", x"FB", x"FF", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"89", x"40", x"40", x"40", x"40", x"60", x"40", x"40", x"89", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"88", x"A8", x"A8", x"88", x"88", x"88", x"88", x"84", x"88", x"D1", x"F5", x"D1", x"F1", x"F5", x"FA", x"FA", x"F5", x"F1", x"D1", x"F5", x"FA", x"FF", x"FF", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"8D", x"40", x"D1", x"F6", x"F6", x"F1", x"84", x"40", x"89", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"B1", x"88", x"88", x"A8", x"68", x"88", x"88", x"A8", x"A8", x"A8", x"D1", x"F5", x"FA", x"FA", x"F5", x"F1", x"D1", x"D1", x"F5", x"D1", x"FA", x"F6", x"D1", x"FB", x"FF", x"D6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"84", x"F5", x"FA", x"FA", x"F9", x"D1", x"64", x"89", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F2", x"E9", x"CD", x"84", x"88", x"88", x"84", x"A8", x"88", x"F1", x"F1", x"F1", x"F6", x"FA", x"FA", x"FA", x"FA", x"F5", x"F1", x"CD", x"CD", x"AD", x"AC", x"D6", x"FA", x"D1", x"F6", x"FA", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F5", x"FA", x"F6", x"F6", x"FA", x"F1", x"D1", x"AD", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F2", x"F2", x"E9", x"E9", x"EE", x"88", x"88", x"88", x"88", x"C8", x"A8", x"D1", x"F5", x"F5", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F5", x"F1", x"F1", x"CC", x"D1", x"F1", x"F6", x"FA", x"F6", x"F6", x"F1", x"F1", x"D1", x"B1", x"D1", x"D1", x"D1", x"D2", x"FF", x"FF", x"D1", x"F6", x"FA", x"FA", x"F5", x"F6", x"FA", x"F5", x"F1", x"CD", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"EE", x"F2", x"EE", x"64", x"88", x"84", x"AD", x"F1", x"AC", x"F5", x"F5", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F1", x"D1", x"F1", x"F6", x"F6", x"FA", x"FA", x"FA", x"F6", x"FA", x"FA", x"F5", x"F1", x"ED", x"F1", x"F1", x"F1", x"F1", x"D1", x"D1", x"F1", x"FA", x"FA", x"FA", x"F5", x"F5", x"FA", x"F6", x"F5", x"D1", x"FB"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"EE", x"EE", x"EE", x"F7", x"D6", x"84", x"88", x"84", x"C9", x"F1", x"F1", x"F1", x"F5", x"FA", x"FA", x"FA", x"FA", x"F6", x"F6", x"F5", x"F1", x"F5", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F6", x"F6", x"F6", x"FA", x"F5", x"F1", x"F1", x"F5", x"F6", x"F6", x"F5", x"F5", x"FA", x"FA", x"FA", x"F6", x"F1", x"F5", x"FA", x"FA", x"F5", x"D1", x"FB"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"A8", x"CD", x"CD", x"CD", x"F1", x"F1", x"F1", x"FA", x"F6", x"F6", x"F6", x"F5", x"F1", x"F1", x"F6", x"FA", x"F5", x"F6", x"F6", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F6", x"F5", x"F6", x"FA", x"F6", x"F1", x"F5", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F6", x"F5", x"F1", x"F1", x"F6", x"F5", x"F5", x"F1", x"FB"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"EE", x"EE", x"CD", x"F2", x"CD", x"88", x"CE", x"F7", x"EE", x"ED", x"F1", x"FA", x"FA", x"F6", x"F5", x"F1", x"F5", x"FA", x"FA", x"FA", x"F6", x"F5", x"F6", x"F6", x"FA", x"FA", x"F6", x"F6", x"F6", x"F6", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F6", x"F5", x"F1", x"F5", x"F1", x"F5", x"F5", x"F6", x"F6", x"F1", x"F1", x"F5", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"F3", x"F2", x"C8", x"B1", x"F7", x"F2", x"ED", x"F5", x"FA", x"FA", x"FA", x"F6", x"F5", x"F6", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F1", x"F5", x"F5", x"F1", x"F1", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F5", x"F6", x"F5", x"F5", x"F6", x"F6", x"F6", x"F6", x"FA", x"F6", x"CD", x"F1", x"D6", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"ED", x"F2", x"EE", x"EE", x"F2", x"F2", x"F7", x"F7", x"EE", x"F2", x"F7", x"F7", x"F2", x"F1", x"FA", x"FA", x"FA", x"F6", x"F5", x"F6", x"F6", x"F6", x"FA", x"FA", x"F5", x"F1", x"F1", x"CD", x"F1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"F5", x"F1", x"F5", x"F1", x"F1", x"F5", x"F6", x"F5", x"F1", x"F1", x"F1", x"F5", x"F1", x"F1", x"F1", x"88", x"D2", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F5", x"ED", x"EE", x"EE", x"EE", x"EE", x"EE", x"D7", x"F7", x"F7", x"EE", x"F7", x"D7", x"F7", x"F2", x"F6", x"FA", x"F6", x"F5", x"F6", x"F6", x"F5", x"F6", x"F6", x"F1", x"F1", x"F1", x"F1", x"CD", x"AC", x"F1", x"F1", x"F5", x"F5", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"AC", x"AD", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"CD", x"D1", x"ED", x"EE", x"EE", x"C9", x"EE", x"F7", x"D7", x"F2", x"EE", x"F2", x"F7", x"D7", x"F2", x"F2", x"F6", x"FA", x"F5", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F5", x"F5", x"F1", x"CD", x"A8", x"AC", x"CD", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"CD", x"CD", x"CD", x"D1", x"F6", x"D6", x"F6", x"FA", x"FA", x"DA", x"D6", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F1", x"F5", x"F1", x"E9", x"ED", x"C9", x"F2", x"F2", x"D7", x"F7", x"F2", x"F2", x"F2", x"F7", x"F7", x"F2", x"D1", x"F5", x"F5", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F5", x"F5", x"F1", x"F1", x"AC", x"88", x"88", x"A8", x"A8", x"A8", x"A8", x"A8", x"A8", x"CC", x"CD", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"F5", x"F1", x"F5", x"ED", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F7", x"D7", x"69", x"44", x"44", x"44", x"B1", x"FA", x"F6", x"F6", x"F6", x"F5", x"F1", x"CD", x"A8", x"64", x"8D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"F1", x"F5", x"F1", x"F5", x"F5", x"CD", x"C9", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F7", x"D7", x"B2", x"24", x"00", x"00", x"24", x"20", x"68", x"D1", x"CD", x"44", x"20", x"20", x"00", x"24", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"CD", x"F1", x"F1", x"F5", x"F5", x"F5", x"ED", x"C5", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F7", x"D7", x"F7", x"8E", x"45", x"00", x"00", x"00", x"00", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B1", x"F5", x"F1", x"F1", x"F1", x"F5", x"F5", x"F1", x"C9", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"8E", x"69", x"69", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"F5", x"F1", x"F1", x"F1", x"F1", x"F1", x"CD", x"EA", x"EE", x"F2", x"F2", x"EE", x"F2", x"CE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"FB", x"D2", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"CD", x"F1", x"ED", x"CC", x"CD", x"AD", x"C9", x"C9", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"CD", x"EE", x"F7", x"F7", x"D2", x"B2", x"89", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"D7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"AD", x"CD", x"AD", x"AD", x"CD", x"C9", x"ED", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"F2", x"EE", x"F2", x"EE", x"EE", x"EE", x"C9", x"C9", x"E9", x"EE", x"EE", x"EE", x"85", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EA", x"EA", x"EE", x"EE", x"EE", x"C9", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"EE", x"C9", x"E9", x"C9", x"EE", x"89", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"CE", x"89", x"64", x"64", x"64", x"65", x"64", x"64", x"A5", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"AD", x"20", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"CE", x"85", x"85", x"85", x"89", x"89", x"89", x"89", x"A5", x"C5", x"E9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"A9", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"C9", x"C9", x"EE", x"EE", x"F2", x"F2", x"F7", x"F7", x"F2", x"CE", x"C5", x"C9", x"EE", x"EE", x"EE", x"F2", x"EE", x"F2", x"EE", x"EE", x"EE", x"E9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"D7", x"F7", x"CE", x"C5", x"C5", x"C9", x"EE", x"CD", x"EE", x"EE", x"EE", x"EE", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"F2", x"EE", x"CE", x"EE", x"EE", x"CD", x"C9", x"C5", x"C5", x"C5", x"C9", x"E9", x"C5", x"C9", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"E9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"F2", x"EE", x"F7", x"D7", x"F2", x"F2", x"EE", x"EA", x"F2", x"C9", x"A5", x"60", x"60", x"C9", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EA", x"EE", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"CE", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"EE", x"ED", x"F2", x"AD", x"00", x"00", x"AD", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F7", x"EE", x"D2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"C9", x"EE", x"AD", x"00", x"00", x"AD", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"EE", x"C9", x"AD", x"00", x"00", x"AD", x"EE", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"C9", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"C9", x"A9", x"00", x"00", x"A9", x"F7", x"F7", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C5", x"C5", x"C9", x"C9", x"E9", x"EE", x"F2", x"F2", x"F3", x"F7", x"D7", x"F7", x"F7", x"D7", x"F7", x"F2", x"CE", x"C5", x"40", x"00", x"00", x"AE", x"F7", x"F3", x"F7", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"C9", x"E9", x"EA", x"F2", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"D7", x"F7", x"D7", x"F7", x"F2", x"E9", x"A0", x"00", x"00", x"00", x"CE", x"F2", x"F2", x"D6", x"F7", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"EE", x"F7", x"D7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"C5", x"A5", x"00", x"00", x"00", x"AD", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"F7", x"D7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"D7", x"F2", x"EE", x"C5", x"A5", x"00", x"00", x"85", x"E9", x"F2", x"F2", x"EE", x"F2", x"F7", x"F7", x"D7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"EE", x"F2", x"F2", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"D7", x"D7", x"F7", x"EE", x"C9", x"C5", x"A5", x"00", x"00", x"85", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F7", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"ED", x"F2", x"F2", x"F2", x"F2", x"F7", x"D7", x"F7", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"D7", x"F2", x"EE", x"C5", x"C5", x"C9", x"65", x"65", x"A9", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F3", x"F7", x"F7", x"F3", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"EE", x"C5", x"C5", x"C5", x"C9", x"E9", x"E9", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F6", x"F7", x"F7", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F2", x"E9", x"C5", x"C9", x"E9", x"E9", x"E9", x"E9", x"CD", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F6", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"F2", x"F6", x"D7", x"D7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"EA", x"C5", x"C5", x"C9", x"C9", x"C9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"EE", x"CE", x"FF", x"D2", x"C5", x"C5", x"C9", x"C9", x"C9", x"E9", x"EA", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"D7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"CE", x"FF", x"FF", x"FF", x"FB", x"C9", x"C5", x"C9", x"E9", x"C9", x"EE", x"CD", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"E9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"D7", x"F7", x"F7", x"D7", x"F7", x"F7", x"D7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"C9", x"C9", x"ED", x"E9", x"EE", x"E9", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"E9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"D7", x"D7", x"F7", x"F7", x"D7", x"D7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"C5", x"C9", x"C9", x"C9", x"C9", x"EA", x"EE", x"CE", x"ED", x"EE", x"EA", x"EA", x"CE", x"EE", x"E9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"D7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C5", x"C5", x"C9", x"E9", x"C9", x"EE", x"EE", x"EE", x"CD", x"CD", x"EE", x"EE", x"EE", x"ED", x"E9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"CD", x"ED", x"EE", x"ED", x"EE", x"E9", x"EE", x"EE", x"EE", x"EE", x"CD", x"EE", x"EE", x"E9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"F2", x"F7", x"F7", x"F3", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"EE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C5", x"C9", x"ED", x"EE", x"EE", x"E9", x"EE", x"EE", x"ED", x"EE", x"EE", x"EE", x"EE", x"EE", x"E9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"F2", x"CE", x"EE", x"EE", x"EE", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"C9", x"CD", x"ED", x"ED", x"EE", x"EE", x"CE", x"ED", x"EE", x"EA", x"EA", x"EE", x"EE", x"E9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EE", x"F2", x"F2", x"F3", x"D7", x"F7", x"F7", x"F7", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"E9", x"EE", x"EE", x"EA", x"CD", x"EE", x"EE", x"EE", x"EE", x"E9", x"E9", x"CE", x"EE", x"E9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"CE", x"EE", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"EE", x"C9", x"C9", x"EE", x"EE", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"EE", x"EE", x"F7", x"D7", x"F7", x"F3", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C9", x"CE", x"EE", x"CE", x"CD", x"EE", x"CE", x"ED", x"EE", x"C9", x"E9", x"E9", x"C9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"CE", x"C5", x"A4", x"CD", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"C9", x"EA", x"EE", x"ED", x"EE", x"EE", x"EE", x"EE", x"E9", x"C9", x"ED", x"EE", x"E9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"A4", x"88", x"A9", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"CE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"EE", x"EA", x"EE", x"E9", x"EE", x"EE", x"E9", x"E9", x"C9", x"EE", x"ED", x"E9", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"A8", x"D1", x"AD", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"C5", x"E9", x"EE", x"E9", x"EA", x"CE", x"EE", x"E9", x"C9", x"C9", x"EE", x"EE", x"C9", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"F1", x"F1", x"CD", x"AD", x"CD", x"CD", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C5", x"ED", x"CD", x"CE", x"EE", x"ED", x"E9", x"C9", x"C9", x"E9", x"EE", x"CE", x"E9", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"D6", x"CD", x"F1", x"F1", x"F1", x"F5", x"F5", x"F1", x"F1", x"F1", x"CD", x"ED", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"C9", x"E9", x"EE", x"EE", x"EE", x"E9", x"C9", x"C9", x"C9", x"E9", x"EE", x"C9", x"E9", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"F6", x"D1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"CD", x"F1", x"F1", x"AD", x"C9", x"C9", x"EE", x"F2", x"F2", x"EE", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"EA", x"E9", x"E9", x"C9", x"C9", x"C9", x"C9", x"CE", x"C9", x"E9", x"F2", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"D2", x"F1", x"F1", x"F5", x"F1", x"F5", x"F5", x"F1", x"D1", x"CD", x"CD", x"D6", x"FF", x"F2", x"C9", x"EE", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"C9", x"C9", x"CD", x"CD", x"A8", x"C9", x"FB", x"FF", x"F7", x"F6", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FB", x"AD", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"CD", x"CD", x"FF", x"FF", x"FF", x"FB", x"C9", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CC", x"CD", x"D1", x"F1", x"CC", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"D6", x"CD", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"F1", x"D1", x"F1", x"ED", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"F6", x"F1", x"F1", x"F5", x"F5", x"F5", x"F1", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"CD", x"CD", x"F1", x"F1", x"F1", x"F1", x"CD", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"CD", x"F1", x"F5", x"F1", x"F5", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"CD", x"F1", x"ED", x"CD", x"ED", x"F1", x"F1", x"F1", x"F1", x"F6", x"FA", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"CD", x"F5", x"F5", x"F5", x"F5", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"D1", x"F1", x"F1", x"ED", x"F1", x"F1", x"D1", x"F1", x"F1", x"F1", x"F1", x"D1", x"D1", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"CD", x"F5", x"F5", x"F5", x"F5", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DF", x"CD", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"D1", x"ED", x"F1", x"ED", x"ED", x"F1", x"ED", x"CD", x"D1", x"D1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FB", x"AD", x"F1", x"F5", x"F5", x"F5", x"F5", x"CD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"A9", x"CD", x"CC", x"CC", x"CC", x"CD", x"CC", x"CD", x"CD", x"CD", x"D1", x"ED", x"F1", x"F1", x"F1", x"ED", x"F1", x"F1", x"F1", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"DA", x"CD", x"F1", x"F5", x"F5", x"F5", x"F5", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"B1", x"B1", x"B1", x"AD", x"B1", x"B1", x"D2", x"D2", x"D1", x"CD", x"CC", x"A8", x"A8", x"AC", x"CD", x"CD", x"AC", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"D1", x"F1", x"F1", x"F5", x"F5", x"D1", x"F1", x"F5", x"F5", x"F1", x"DA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DA", x"D6", x"DA", x"FA", x"DB", x"DA", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"D1", x"D1", x"D1", x"D1", x"CD", x"AC", x"AC", x"CD", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
);
constant PinkPunch_bmp: PinkPunch_bmp_array := (
("0000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000001111100000"),
("0000000000000000000000000000000000000000001111111000000000000111111110000"),
("0000000000000000000000000000000000000000111111111100000000001111111111000"),
("0000000000000000000000000000000000000001111111111110000000001111111111000"),
("0000000000000000000000000000000000000001111111111111000000001111111111100"),
("0000000000000000000000000000000000000011111111111111100000001111111111100"),
("0000000000000000000000000000000000000011111111111111110000001111111111110"),
("0000000000000000000000000000000000000011111111111111110000001111111111110"),
("0000000000000000000000000000000011111111111111111111011000000111111111110"),
("0000000000000000000000000000000111111111111111111111011000000001111111110"),
("0000000000000000000000000000011111111111111111111110010000000001111111110"),
("0000000000000000000000000011111111111111111111111110110000000001111111110"),
("0000000000000000000000011111111111111111111111111111100000000001111111110"),
("0000000000000000000011111111111111111111111111111111111111110011111111110"),
("0000000000000000000011111111111111111111111111111111111111111111111111111"),
("0000000000000000000111111111111111111111111111111111111111111111111111111"),
("0000000000000000000111111111111111111111111111111111111111111111111111111"),
("0000000000000000000111111111111111111111111111111111111111111111111111110"),
("0000000000000000000111111111111111111111111111111111111111111111111111110"),
("0000000000000000001111111111111111111111111111111111111111111111111111100"),
("0000000000000000001111111111111111111111111111111111111111111111111111000"),
("0000000000000000011111111111111111111111111111111111111111111111111110000"),
("0000000000000000011111111111111111111111111111111111111111100000000000000"),
("0000000000000000111111111111111111111111111111111100000000000000000000000"),
("0000000000000000111111111111111111111111111111111110000000000000000000000"),
("0000000000000001111111111111111111111111111111111111000000000000000000000"),
("0000000000000001111111111111111111111111111111111111100000000000000000000"),
("0000000000000001111111111111111111111111111111111111110000000000000000000"),
("0000000000000000111111111111111111111111111111111111110000000000000000000"),
("0000000000000000011111111111111111111111111111111111100000000000000000000"),
("0000000000000000000000000111111111111111111111111111100000000000000000000"),
("0000000000000000000000000111111111111111111111111110000000000000000000000"),
("0000000000000000000000000111111111111111111111111100000000000000000000000"),
("0000000000000000000000000111111111111111111111111000000000000000000000000"),
("0000000000000000000000001111111111111111111111110000000000000000000000000"),
("0000000000000000000000011111111111111111111111100000000000000000000000000"),
("0000000000000000000000111111111111111111111111000000000000000000000000000"),
("0000000000000000000001111111111111111111111111000000000000000000000000000"),
("0000000000000000000001111111111111111111111111100000000000000000000000000"),
("0000000000000000000001111111111111111111111111110000000000000000000000000"),
("0000000000000000000000111111111111111111111111111000000000000000000000000"),
("0000000000000000000000011111111111111111111111111000000000000000000000000"),
("0000000000000000000000011111111111111111111111111100000000000000000000000"),
("0000000000000000000000111111111111111111111111111110000000000000000000000"),
("0000000000000000000001111111111111111111111111111111000000000000000000000"),
("0000000000000000000011111111111111111111111111111111100000000000000000000"),
("0000000000000000000111111111111111111111111111111111110000000000000000000"),
("0000000000000000000111111111111111111111111111111111111000000000000000000"),
("0000000000000000000111111111111111111111111111111111111100000000000000000"),
("0000000000000000000111111111111111111111111111111111111100000000000000000"),
("0000000000000000001111111111111111110111111111111111111110000000000000000"),
("0000000000000000011111111111111111100011111111111111111110000000000000000"),
("0000000000000000111111111111111111000000111111111111111110000000000000000"),
("0000000000000011111111111111111110000000011111111111111110000000000000000"),
("0000000000000011111111111111111100000000001111111111111110000000000000000"),
("0000000000000111111111111111111000000000011111111111111110000000000000000"),
("0000000000001111111111111111111000000000011111111111111110000000000000000"),
("0000000000011111111111111111100000000000001111111111111110000000000000000"),
("0000000000111111111111111111000000000000001111111111111110000000000000000"),
("0000000011111111111111111110000000000000001111111111111110000000000000000"),
("0000000111111111111111111100000000000000001111111111111110000000000000000"),
("0000001111111111111111111000000000000000001111111111111110000000000000000"),
("0000001111111111111111110000000000000000001111111111111110000000000000000"),
("0000000111111111111111100000000000000000001111111111111110000000000000000"),
("0000001111111111111111000000000000000000001111111111111110000000000000000"),
("0011111111111111111110000000000000000000001111111111111110000000000000000"),
("0111111111111111111100000000000000000000000111111111111110000000000000000"),
("0111111111111011111000000000000000000000000011111111011010000000000000000"),
("0111111111110001110000000000000000000000000011111110000000000000000000000"),
("0011111111110000000000000000000000000000000011111110000000000000000000000"),
("0001111111100000000000000000000000000000000111111111100000000000000000000"),
("0000111111100000000000000000000000000000001111111111111000000000000000000"),
("0000111111000000000000000000000000000000011111111111111110000000000000000"),
("0000111111000000000000000000000000000000111111111111111111110000000000000"),
("0011111111100000000000000000000000000000011111111111111111111100000000000"),
("0011111111100000000000000000000000000000001111111111111111111100000000000"),
("0001111111111100000000000000000000000000000000000000111111111000000000000"),
("0000111111111000000000000000000000000000000000000000000000000000000000000")
);
constant PinkShoot_X_size : integer := 90;
constant PinkShoot_Y_size : integer := 83;
type PinkShoot_color_array is array(0 to PinkShoot_Y_size - 1 , 0 to PinkShoot_X_size - 1) of std_logic_vector(7 downto 0);
type PinkShoot_bmp_array is array(0 to PinkShoot_Y_size - 1 , 0 to PinkShoot_X_size - 1) of std_logic;
constant PinkShoot_colors: PinkShoot_color_array := (
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AD", x"88", x"88", x"88", x"88", x"84", x"88", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"88", x"88", x"88", x"88", x"88", x"84", x"88", x"88", x"88", x"8C", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"84", x"84", x"88", x"88", x"84", x"88", x"88", x"88", x"84", x"88", x"88", x"88", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"DA", x"FF", x"FF", x"F1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"88", x"88", x"88", x"88", x"88", x"CD", x"AC", x"AC", x"AC", x"88", x"88", x"64", x"B1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F5", x"D1", x"D6", x"FF", x"F5", x"F5", x"FA", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AC", x"88", x"88", x"88", x"A8", x"A8", x"D1", x"D1", x"44", x"B5", x"F5", x"AC", x"88", x"AD", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"D5", x"D2", x"F6", x"F5", x"F2", x"D6", x"FA", x"FA", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"88", x"88", x"CC", x"8C", x"84", x"A8", x"D1", x"8D", x"00", x"68", x"F6", x"F1", x"CC", x"FB", x"D6", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F5", x"D1", x"88", x"64", x"89", x"D1", x"AC", x"D5", x"F1", x"D1", x"FB", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"AD", x"AD", x"AD", x"AC", x"88", x"A4", x"CC", x"F6", x"F5", x"AC", x"F1", x"F5", x"D1", x"44", x"00", x"D1", x"FA", x"D1", x"F6", x"FF", x"8C", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"F5", x"AD", x"64", x"40", x"40", x"40", x"64", x"64", x"F5", x"D5", x"D6", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"88", x"A8", x"88", x"A8", x"88", x"88", x"88", x"A9", x"88", x"D1", x"F5", x"D5", x"F6", x"F6", x"F6", x"AD", x"24", x"44", x"F1", x"FA", x"FF", x"FF", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"D1", x"D1", x"64", x"40", x"60", x"60", x"60", x"40", x"40", x"88", x"F1", x"F1", x"F6", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DA", x"88", x"88", x"AC", x"A8", x"88", x"88", x"88", x"84", x"84", x"88", x"D1", x"D1", x"D1", x"F1", x"F5", x"FA", x"F6", x"F5", x"F1", x"D1", x"F5", x"FB", x"FB", x"DA", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"88", x"40", x"20", x"40", x"40", x"40", x"40", x"60", x"60", x"60", x"89", x"D1", x"D2", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"DB", x"88", x"88", x"A8", x"A8", x"88", x"88", x"A9", x"A9", x"AD", x"AD", x"EE", x"F2", x"D2", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F6", x"FA", x"F6", x"CE", x"A4", x"F2", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"FA", x"FA", x"FA", x"FB", x"FF", x"D6", x"A8", x"88", x"64", x"40", x"40", x"40", x"40", x"40", x"60", x"40", x"40", x"D1", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"F2", x"EE", x"EA", x"A9", x"84", x"88", x"88", x"88", x"88", x"AD", x"F7", x"F3", x"F2", x"F2", x"F2", x"F2", x"F3", x"F7", x"F7", x"F2", x"F2", x"F2", x"D2", x"D2", x"F7", x"D2", x"69", x"65", x"89", x"C9", x"C5", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"FA", x"F6", x"F5", x"F5", x"F1", x"F1", x"F5", x"F6", x"FA", x"FA", x"F6", x"F6", x"F5", x"88", x"40", x"60", x"40", x"40", x"40", x"20", x"8D", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"F6", x"EE", x"C9", x"EE", x"CD", x"88", x"88", x"88", x"88", x"AD", x"AD", x"F7", x"F7", x"F7", x"F7", x"D6", x"F7", x"D7", x"F7", x"F7", x"F3", x"F7", x"F7", x"F7", x"F7", x"F2", x"CE", x"44", x"44", x"8D", x"CD", x"CD", x"CD", x"C9", x"F1", x"F6", x"F5", x"D5", x"D5", x"D1", x"FB", x"FF", x"F6", x"F6", x"F6", x"FA", x"F6", x"F6", x"F6", x"F6", x"FA", x"FA", x"F5", x"F6", x"F6", x"F6", x"FA", x"B1", x"40", x"60", x"40", x"40", x"40", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"EE", x"EE", x"EE", x"F2", x"CD", x"84", x"88", x"88", x"F6", x"B2", x"CD", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F7", x"F7", x"D7", x"D7", x"F6", x"D2", x"44", x"44", x"D6", x"FA", x"F6", x"F6", x"F5", x"F1", x"F1", x"F1", x"F1", x"F5", x"F1", x"F1", x"D1", x"F6", x"FA", x"FA", x"FA", x"F6", x"F6", x"F6", x"FA", x"FA", x"FA", x"F6", x"FA", x"F6", x"FA", x"FA", x"F5", x"CC", x"40", x"40", x"40", x"44", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"EE", x"F2", x"F7", x"AD", x"84", x"88", x"88", x"F7", x"D7", x"D7", x"F7", x"D7", x"F7", x"D7", x"D7", x"F7", x"F7", x"F2", x"F7", x"F7", x"F7", x"F2", x"EE", x"A9", x"20", x"00", x"D6", x"F6", x"F6", x"F6", x"F6", x"FA", x"F5", x"D1", x"F1", x"F6", x"F6", x"F6", x"F6", x"FA", x"F6", x"F6", x"F6", x"F5", x"F6", x"FA", x"FA", x"FA", x"FA", x"FA", x"F6", x"F6", x"F1", x"F1", x"F1", x"CD", x"84", x"40", x"40", x"89", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"F2", x"EE", x"EE", x"EE", x"F2", x"D2", x"88", x"D1", x"AD", x"D2", x"D6", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F6", x"F2", x"F2", x"F2", x"F2", x"F2", x"CE", x"89", x"89", x"24", x"44", x"F1", x"F1", x"F5", x"F5", x"F6", x"F6", x"FA", x"F5", x"F1", x"F5", x"F5", x"F5", x"F6", x"F6", x"F6", x"F1", x"F1", x"F1", x"F5", x"F6", x"F5", x"F6", x"F5", x"F5", x"F5", x"F1", x"F1", x"CD", x"A8", x"D1", x"8D", x"B1", x"B2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F7", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"AD", x"A8", x"D2", x"D2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F3", x"F3", x"F2", x"F3", x"F6", x"F7", x"F7", x"F7", x"F2", x"44", x"00", x"00", x"B1", x"F5", x"F1", x"F6", x"FA", x"FA", x"FA", x"FA", x"F6", x"FA", x"FA", x"F6", x"F6", x"F5", x"F6", x"F6", x"F5", x"F5", x"F6", x"F5", x"F6", x"F5", x"F1", x"F1", x"F1", x"F1", x"CD", x"AC", x"B1", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"88", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"CE", x"64", x"00", x"D1", x"F1", x"F6", x"FA", x"FA", x"F6", x"F6", x"FA", x"FA", x"FA", x"F6", x"F6", x"F6", x"F6", x"FA", x"F6", x"FA", x"FA", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"CC", x"AD", x"DA", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D1", x"F1", x"F2", x"EE", x"EE", x"F2", x"F2", x"DB", x"F2", x"F2", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F2", x"AE", x"20", x"00", x"89", x"F1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"F1", x"F1", x"AD", x"CC", x"CD", x"AD", x"AD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F1", x"ED", x"EE", x"EE", x"EE", x"CE", x"F2", x"D7", x"F7", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"44", x"00", x"00", x"8D", x"F1", x"F1", x"F1", x"F5", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"CD", x"CD", x"CD", x"CD", x"CC", x"CD", x"F1", x"B1", x"D1", x"AD", x"8D", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"D1", x"ED", x"EE", x"EE", x"E9", x"E9", x"F2", x"F7", x"F7", x"F2", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F3", x"F7", x"D7", x"D2", x"45", x"00", x"88", x"CD", x"CD", x"CD", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"ED", x"CD", x"D1", x"D1", x"D6", x"D6", x"D6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"F1", x"F5", x"F5", x"ED", x"CA", x"C9", x"EE", x"F2", x"F7", x"F7", x"F7", x"F2", x"F2", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F3", x"F7", x"F7", x"D2", x"44", x"00", x"88", x"F1", x"CC", x"CD", x"CD", x"A8", x"A8", x"A8", x"A8", x"AC", x"CC", x"D1", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"F1", x"F1", x"F5", x"F1", x"CD", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F3", x"D7", x"D7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F7", x"CD", x"00", x"00", x"24", x"AD", x"ED", x"AD", x"44", x"84", x"C5", x"A9", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"CD", x"F1", x"F5", x"F5", x"F1", x"F1", x"C9", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F6", x"EE", x"F3", x"F2", x"89", x"20", x"00", x"00", x"24", x"24", x"64", x"C9", x"C5", x"C9", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"D1", x"F1", x"F1", x"F1", x"F5", x"F5", x"C9", x"E9", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"F7", x"D2", x"CA", x"64", x"40", x"40", x"C5", x"C5", x"C9", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"F6", x"F1", x"F1", x"F5", x"F5", x"F5", x"ED", x"C9", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"D2", x"CE", x"D2", x"F2", x"ED", x"EA", x"C9", x"E9", x"C5", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"F1", x"C9", x"EE", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EA", x"CD", x"CE", x"C9", x"C9", x"C9", x"C9", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"CD", x"D0", x"CD", x"CC", x"AC", x"AD", x"C5", x"C9", x"EE", x"EE", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"C9", x"C9", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"AD", x"CD", x"AD", x"AD", x"CD", x"C9", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"EE", x"EE", x"EA", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"EE", x"EA", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"AD", x"65", x"64", x"84", x"64", x"64", x"84", x"65", x"69", x"A9", x"EE", x"EE", x"EE", x"EE", x"A9", x"89", x"89", x"64", x"85", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"AD", x"84", x"64", x"89", x"89", x"89", x"89", x"85", x"64", x"60", x"44", x"64", x"64", x"60", x"20", x"00", x"00", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"CE", x"E9", x"E9", x"EE", x"F2", x"F2", x"F3", x"F7", x"F7", x"F2", x"CE", x"AD", x"A9", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"F2", x"F7", x"F7", x"F7", x"F3", x"F7", x"F7", x"F2", x"CE", x"CE", x"CE", x"44", x"00", x"CE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"F2", x"EE", x"F2", x"F2", x"EE", x"F2", x"F7", x"D7", x"F2", x"EE", x"CE", x"EE", x"C9", x"EE", x"F2", x"F2", x"F2", x"69", x"00", x"CE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"E9", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"D6", x"EE", x"F2", x"D7", x"F7", x"F3", x"F2", x"EE", x"EE", x"EE", x"F2", x"65", x"00", x"85", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"EE", x"EE", x"F2", x"65", x"00", x"24", x"EE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"EE", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F2", x"C9", x"F2", x"65", x"00", x"20", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"D2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"E9", x"EE", x"69", x"00", x"20", x"EE", x"CE", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"EE", x"EE", x"F2", x"F2", x"D2", x"EE", x"F2", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"E9", x"E9", x"65", x"00", x"20", x"CE", x"D7", x"F7", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"C5", x"C5", x"E9", x"C9", x"E9", x"EE", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F2", x"C9", x"A5", x"20", x"00", x"24", x"F2", x"F3", x"F7", x"F7", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"E9", x"C9", x"E9", x"CE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F6", x"EE", x"E9", x"60", x"00", x"00", x"24", x"F2", x"F2", x"F2", x"F7", x"D7", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"CD", x"EE", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F2", x"EE", x"C5", x"64", x"00", x"00", x"44", x"F2", x"F2", x"F2", x"F2", x"F7", x"D7", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F6", x"CD", x"EE", x"F2", x"F6", x"F7", x"F3", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"EE", x"E9", x"C5", x"64", x"00", x"00", x"A9", x"EE", x"EE", x"F2", x"EE", x"F2", x"F7", x"F7", x"F2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"EE", x"EE", x"EE", x"EE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"EE", x"A5", x"C9", x"64", x"00", x"00", x"C9", x"EE", x"F2", x"F2", x"F2", x"F2", x"F3", x"D7", x"D7", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"EE", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"D7", x"F7", x"F7", x"F7", x"F2", x"C9", x"C5", x"C9", x"A9", x"64", x"65", x"CE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F6", x"F3", x"F3", x"F7", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"EE", x"F2", x"F6", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F2", x"EE", x"C5", x"C5", x"C9", x"E9", x"E9", x"E9", x"EA", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F3", x"F7", x"F2", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CA", x"EE", x"F2", x"F2", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"C9", x"C5", x"C9", x"E9", x"C9", x"E9", x"C9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F6", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"EE", x"F2", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F2", x"C9", x"C5", x"C5", x"C9", x"C9", x"E9", x"ED", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"F2", x"EE", x"EE", x"F2", x"F2", x"D2", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F2", x"CA", x"D6", x"F6", x"C5", x"C5", x"C9", x"C9", x"E9", x"E9", x"E9", x"CE", x"EE", x"EA", x"EE", x"EE", x"CD", x"CE", x"CE", x"EE", x"F2", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"D7", x"D7", x"F7", x"D7", x"F7", x"CA", x"F6", x"FF", x"FF", x"FB", x"CE", x"C5", x"C9", x"C9", x"C9", x"C9", x"EE", x"EE", x"EE", x"CE", x"EA", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"E9", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"C5", x"C9", x"C9", x"EE", x"EA", x"EE", x"C9", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"CD", x"EE", x"EE", x"CA", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"D7", x"F7", x"F7", x"D7", x"F2", x"F2", x"F2", x"F2", x"C9", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"C9", x"C9", x"C9", x"C9", x"C9", x"EE", x"EE", x"EE", x"CE", x"EE", x"ED", x"EE", x"EE", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EA", x"F2", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F7", x"F3", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"C5", x"C9", x"C9", x"E9", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"EE", x"EE", x"F2", x"F2", x"F2", x"D7", x"F7", x"F7", x"F7", x"F2", x"F2", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"C9", x"E9", x"EE", x"ED", x"EE", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"EE", x"EE", x"F2", x"F7", x"F7", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"E9", x"E9", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"C9", x"C9", x"C9", x"EE", x"E9", x"EE", x"CE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"EE", x"EE", x"C9", x"F2", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"C9", x"EE", x"CD", x"EE", x"EE", x"EE", x"EE", x"EE", x"E9", x"EE", x"ED", x"EE", x"CE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CE", x"EE", x"F2", x"F2", x"D7", x"D7", x"F7", x"F7", x"F6", x"F2", x"F2", x"F2", x"EE", x"EE", x"F2", x"EE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EA", x"EE", x"EE", x"EE", x"EE", x"E9", x"EE", x"CE", x"EE", x"C9", x"E9", x"EA", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EE", x"F2", x"F2", x"F7", x"D7", x"F7", x"F7", x"F7", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"E9", x"EE", x"E9", x"EE", x"EE", x"EE", x"EE", x"CE", x"EE", x"C9", x"EA", x"EE", x"CE", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"F2", x"EE", x"EE", x"F2", x"F7", x"F7", x"F7", x"F3", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"EE", x"EA", x"C9", x"EE", x"CD", x"EE", x"EE", x"EE", x"ED", x"E9", x"C9", x"EA", x"EE", x"C9", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"C5", x"A9", x"ED", x"F2", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"F2", x"CE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CE", x"E9", x"EE", x"ED", x"EE", x"CE", x"EE", x"CE", x"EE", x"C9", x"CA", x"EE", x"EE", x"CD", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"A4", x"A8", x"AD", x"EE", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F2", x"EE", x"EE", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"C9", x"ED", x"E9", x"EE", x"CE", x"CD", x"EE", x"EA", x"C9", x"E9", x"ED", x"EE", x"EE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"CD", x"CD", x"CD", x"EE", x"EE", x"EE", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"CA", x"EE", x"EE", x"EE", x"EE", x"CE", x"ED", x"C9", x"C9", x"C9", x"C9", x"EE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D6", x"CD", x"F1", x"CD", x"CD", x"CD", x"CD", x"CD", x"F2", x"EE", x"F2", x"F2", x"F2", x"F2", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"C9", x"E9", x"EA", x"EE", x"EE", x"EA", x"C9", x"C9", x"C9", x"E9", x"EE", x"CE", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"D2", x"CD", x"F1", x"F1", x"F1", x"F5", x"F1", x"F1", x"F1", x"F1", x"CD", x"ED", x"EE", x"F2", x"F2", x"F2", x"EE", x"EE", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"D2", x"E9", x"ED", x"EE", x"CD", x"CE", x"C9", x"C5", x"C5", x"C9", x"C9", x"CD", x"ED", x"CE", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"D2", x"F1", x"F1", x"F5", x"F5", x"F5", x"F1", x"D1", x"D1", x"F5", x"D1", x"CD", x"C9", x"C9", x"F2", x"F2", x"F2", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"F2", x"CA", x"EE", x"EA", x"E9", x"A9", x"C9", x"C5", x"CD", x"CD", x"E9", x"ED", x"F2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"CD", x"F1", x"F5", x"F5", x"F1", x"F1", x"F5", x"F1", x"CD", x"CD", x"CD", x"DA", x"FB", x"C9", x"C9", x"EE", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"C9", x"C9", x"AD", x"CD", x"CD", x"A8", x"CE", x"FB", x"FB", x"C9", x"CE", x"FF", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"D6", x"D1", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"F1", x"CD", x"D6", x"FF", x"FF", x"FB", x"C9", x"EE", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"AD", x"CD", x"CD", x"F1", x"D1", x"AD", x"D2", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"DB", x"CD", x"F1", x"F5", x"F5", x"F5", x"F1", x"F5", x"F5", x"CD", x"D6", x"FF", x"FF", x"FF", x"FF", x"F7", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"F1", x"F1", x"F1", x"D1", x"CD", x"D2", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"F6", x"CD", x"F1", x"F5", x"F6", x"F5", x"F5", x"F1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"CD", x"CD", x"CD", x"F1", x"ED", x"F1", x"D1", x"CD", x"D6", x"FB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"CD", x"F1", x"F5", x"F1", x"F5", x"F1", x"CD", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"F1", x"F1", x"ED", x"D1", x"D1", x"F1", x"F1", x"F1", x"F1", x"D1", x"D1", x"F6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"D1", x"F1", x"F5", x"F5", x"F5", x"F1", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"CD", x"ED", x"D1", x"ED", x"ED", x"D1", x"F1", x"ED", x"D1", x"D1", x"F1", x"F1", x"F1", x"D1", x"D1", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"D1", x"F1", x"F5", x"F5", x"F1", x"F5", x"D1", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"CD", x"ED", x"D1", x"F1", x"F1", x"F1", x"F1", x"ED", x"F1", x"F1", x"D1", x"F1", x"F1", x"F1", x"CD", x"CD", x"D1", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"D1", x"F1", x"F5", x"F6", x"F5", x"F1", x"CD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FA", x"AC", x"CC", x"CC", x"CD", x"CC", x"CC", x"CC", x"CD", x"CD", x"CD", x"ED", x"F1", x"ED", x"F1", x"D1", x"ED", x"F1", x"F5", x"CD", x"AD", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"F1", x"F5", x"F5", x"F5", x"F5", x"F5", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B1", x"AD", x"AD", x"AD", x"AD", x"AD", x"D1", x"D6", x"D1", x"CD", x"CD", x"CD", x"CD", x"AD", x"D1", x"F1", x"D1", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"D1", x"F1", x"F5", x"F5", x"F1", x"D1", x"F5", x"F5", x"F6", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FB", x"FB", x"FB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FB", x"CD", x"CD", x"CD", x"CD", x"CD", x"AD", x"AD", x"D1", x"D6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF"),
( x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF")
);
constant PinkShoot_bmp: PinkShoot_bmp_array := (
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000111111111111100000000000000000000000000011001100000"),
("000000000000000000000000000000000000001111111111111100000000000000000000000000111011100000"),
("000000000000000000000000000000000000001111111111111110000000000000000000000000111111111000"),
("000000000000000000000000000000000000011111111111111111000000000000000000000011111111111100"),
("000000000000000000000000000000001111111111111111111101000000000000000000000111111111111000"),
("000000000000000000000000000000111111111111111111111001000000000000000000001111111111111100"),
("000000000000000000000000000011111111111111111111111111000000000000000000001111111111111100"),
("000000000000000000000000011111111111111111111111111111100000000000111111101111111111111000"),
("000000000000000000000011111111111111111111111111111111110000000011111111111111111111110000"),
("000000000000000000001111111111111111111111111111111111111111110111111111111111111111100000"),
("000000000000000000001111111111111111111111111111111111111111111111111111111111111111000000"),
("000000000000000000011111111111111111111111111111111111111111111111111111111111111100000000"),
("000000000000000000111111111111111111111111111111111111111111111111111111111111111000000000"),
("000000000000000000111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000000000011111111111111111111111111111111111111111111111111111111100000000000000"),
("000000000000000000111111111111111111111111111111111111111111111111111111100000000000000000"),
("000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000"),
("000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000"),
("000000000000000011111111111111111111111111111111111111111110000000000000000000000000000000"),
("000000000000000111111111111111111111111111111111111111110000000000000000000000000000000000"),
("000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000"),
("000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000"),
("000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000"),
("000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000"),
("000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000"),
("000000000000000001111111111111111111111111111110000000000000000000000000000000000000000000"),
("000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000"),
("000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000"),
("000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000"),
("000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000"),
("000000000000000000000001111111111111111111111000000000000000000000000000000000000000000000"),
("000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000"),
("000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000"),
("000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000"),
("000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000"),
("000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000"),
("000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000"),
("000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000"),
("000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000"),
("000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000"),
("000000000000000000001111111111111111111111111111111110000000000000000000000000000000000000"),
("000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000"),
("000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000"),
("000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000"),
("000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000"),
("000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000"),
("000000000000000001111111111111111111111111111111111111111000000000000000000000000000000000"),
("000000000000000011111111111111111110011111111111111111111000000000000000000000000000000000"),
("000000000000000111111111111111111100000111111111111111111000000000000000000000000000000000"),
("000000000000001111111111111111111000000011111111111111111000000000000000000000000000000000"),
("000000000000011111111111111111111000000001111111111111111000000000000000000000000000000000"),
("000000000000111111111111111111110000000011111111111111111000000000000000000000000000000000"),
("000000000001111111111111111111100000000011111111111111111000000000000000000000000000000000"),
("000000000011111111111111111111000000000000111111111111111000000000000000000000000000000000"),
("000000000111111111111111111100000000000000111111111111111000000000000000000000000000000000"),
("000000001111111111111111111000000000000000111111111111111000000000000000000000000000000000"),
("000000111111111111111111110000000000000000111111111111111000000000000000000000000000000000"),
("000000111111111111111111100000000000000000111111111111111000000000000000000000000000000000"),
("000000111111111111111111000000000000000000111111111111110000000000000000000000000000000000"),
("000000011111111111111110000000000000000000111111111111110000000000000000000000000000000000"),
("000000111111111111111100000000000000000000111111111111110000000000000000000000000000000000"),
("001111111111111111111000000000000000000000111111111111110000000000000000000000000000000000"),
("011111111111111111110000000000000000000000011111111111110000000000000000000000000000000000"),
("011111111111111111100000000000000000000000001111111111101000000000000000000000000000000000"),
("011111111111001111000000000000000000000000001111111000000000000000000000000000000000000000"),
("011111111111000010000000000000000000000000001111111100000000000000000000000000000000000000"),
("001111111110000000000000000000000000000000111111111111000000000000000000000000000000000000"),
("000111111110000000000000000000000000000001111111111111100000000000000000000000000000000000"),
("000111111100000000000000000000000000000001111111111111111000000000000000000000000000000000"),
("000111111100000000000000000000000000000011111111111111111111000000000000000000000000000000"),
("000111111100000000000000000000000000000011111111111111111111100000000000000000000000000000"),
("000111111110000000000000000000000000000001111111111111111111100000000000000000000000000000"),
("000111111111100000000000000000000000000000000000000111100000000000000000000000000000000000"),
("000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);

begin
process ( RESETn, CLK)

  	variable current_color : std_logic_vector(7 downto 0);
	variable pixel_valid : std_logic;
	
	variable bCoord_X : integer := 0;-- offset from start position 
	variable bCoord_Y : integer := 0;

	variable drawing_X : std_logic := '0';
	variable drawing_Y : std_logic := '0';

	--		
	variable objectEndX : integer;
	variable objectEndY : integer;

   begin
	if RESETn = '0' then
	   mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;
		pixel_valid := '0';

	elsif rising_edge(CLK) then
	
		if(is_game_over = '1' and player_won = '1') then 
			objectEndX	:= 	ObjectStartX + PinkWon_X_size;
		elsif(is_game_over = '1' ) then 
			objectEndX	:= 	ObjectStartX + PinkDead_X_size;
		elsif(PlayerState = player_state_idle or PlayerState = player_state_move_left or PlayerState = player_state_move_right) then 
				objectEndX	:= 	ObjectStartX + PinkIdle_X_size;
		elsif(PlayerState = player_state_kick) then
				objectEndX := ObjectStartX + PinkKick_X_size;
		elsif(PlayerState = player_state_duck) then 
				objectEndX := ObjectStartX + PinkDucking_X_size;
		elsif(PlayerState = player_state_punch) then 
				objectEndX := ObjectStartX + PinkPunch_X_size;	
		else -- PlayerState = player_state_shoot
				objectEndX := ObjectStartX + PinkShoot_X_size;
		end if;
		
		if(is_game_over = '1' and player_won = '1') then 
			objectEndY	:= 	ObjectStartY + PinkWon_Y_size;
		elsif(is_game_over = '1') then 
			objectEndY	:= 	ObjectStartY + PinkDead_Y_size;
		elsif(PlayerState = player_state_idle or PlayerState = player_state_move_left or PlayerState = player_state_move_right) then 
				objectEndY	:= 	ObjectStartY + PinkIdle_Y_size;
		elsif(PlayerState = player_state_kick) then
				objectEndY := ObjectStartY + PinkKick_Y_size;
		elsif(PlayerState = player_state_duck) then 
				objectEndY := ObjectStartY + PinkDucking_Y_size;
		elsif(PlayerState = player_state_punch) then 
				objectEndY := ObjectStartY + PinkPunch_Y_size;	
		else -- PlayerState = player_state_shoot
				objectEndY := ObjectStartY + PinkShoot_Y_size;
		end if;
	
		if((oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX)) then
			drawing_X	:= '1';
		else 
			drawing_X	:= '0';
		end if;
		
		if((oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY)) then 
			drawing_Y	:= '1';
		else 
			drawing_Y	:= '0';
		end if;

		if(drawing_X = '1' and  drawing_Y = '1' and player_direction = player_direction_right_to_left) then
			bCoord_X 	:= (ObjectEndX - oCoord_X);
		elsif(drawing_X = '1' and  drawing_Y = '1') then 
			bCoord_X 	:= (oCoord_X - ObjectStartX);
		else
			bCoord_X 	:= 0;
		end if;
		
		if( drawing_X = '1' and  drawing_Y = '1') then 
			bCoord_Y 	:= (oCoord_Y - ObjectStartY);
		else
			bCoord_Y 	:= 0;
		end if;
		
		if(is_game_over = '1' and player_won = '1') then 
			current_color := PinkWon_colors(bCoord_Y , bCoord_X);
			pixel_valid := PinkWon_bmp(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
		elsif(is_game_over = '1' ) then 
			current_color := PinkDead_colors(bCoord_Y , bCoord_X);
			pixel_valid := PinkDead_bmp(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
		else
			case PlayerState is
				when  player_state_idle | player_state_move_left | player_state_move_right =>
					--current_color := X"66"; -- yellow
					current_color := PinkIdle_colors(bCoord_Y , bCoord_X);
					pixel_valid := PinkIdle_bmp(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
				when player_state_duck =>
					--current_color := X"E0"; -- red
					current_color := PinkDucking_colors(bCoord_Y , bCoord_X);
					pixel_valid := PinkDucking_bmp(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
				when player_state_shoot =>
					--current_color := X"07";
					--shoot_colors
					current_color := PinkShoot_colors(bCoord_Y , bCoord_X);
					pixel_valid := PinkShoot_bmp(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
				when player_state_punch =>
					current_color := PinkPunch_colors(bCoord_Y , bCoord_X);
					pixel_valid := PinkPunch_bmp(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
				when player_state_kick =>
					current_color := PinkKick_colors(bCoord_Y , bCoord_X);
					pixel_valid := PinkKick_bmp(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
				when others =>
					current_color := X"FF";
					pixel_valid := '0';
			end case;
		end if;
			
		mVGA_RGB				<=  current_color;	--get from colors table 
		drawing_request	<=  pixel_valid; -- get from mask table if inside rectangle  
	end if;

  end process;

		
end behav;		
		
