library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;

package MAIN_MENU_PCKG is 

constant press_S_X_size : integer := 250;
constant press_S_Y_size : integer := 25;
type press_S_color_array is array(0 to press_S_Y_size - 1 , 0 to press_S_X_size - 1) of std_logic_vector(7 downto 0);
constant press_S_colors: press_S_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00"),
( x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"24", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"24", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"24", x"24", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"24", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"24", x"24", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"24", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"24", x"24", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"24", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"24", x"49", x"49", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"00", x"00", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"49", x"24", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"24", x"24", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"49", x"24", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"24", x"49", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"24", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"24", x"24", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"24", x"24", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"24", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);



constant OPTIONS_X_size : integer := 139;
constant OPTIONS_Y_size : integer := 35;
type OPTIONS_color_array is array(0 to OPTIONS_Y_size - 1 , 0 to OPTIONS_X_size - 1) of std_logic_vector(7 downto 0);
constant OPTIONS_colors: OPTIONS_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"75", x"75", x"71", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"71", x"00", x"00", x"00", x"00", x"00", x"24", x"71", x"4D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"71", x"71", x"71", x"4D", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"72", x"49", x"00", x"00", x"00", x"24", x"71", x"4D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"71", x"24", x"00", x"00", x"00", x"00", x"24", x"71", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"71", x"75", x"71", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"28", x"71", x"71", x"71", x"75", x"76", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"72", x"71", x"71", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"00", x"00", x"00", x"00", x"24", x"71", x"6D", x"00", x"00"),
( x"00", x"00", x"00", x"24", x"4D", x"76", x"5D", x"3D", x"3D", x"3D", x"7A", x"49", x"00", x"00", x"00", x"00", x"44", x"71", x"76", x"00", x"00", x"24", x"7A", x"5D", x"28", x"00", x"00", x"00", x"49", x"7A", x"3D", x"71", x"00", x"00", x"00", x"00", x"00", x"48", x"71", x"59", x"3D", x"3D", x"3D", x"5D", x"75", x"24", x"00", x"00", x"00", x"6D", x"5A", x"3D", x"71", x"00", x"24", x"4D", x"7A", x"3D", x"76", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"5A", x"3D", x"7A", x"71", x"24", x"24", x"4D", x"76", x"3D", x"76", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"75", x"5D", x"3D", x"5D", x"76", x"24", x"00", x"00", x"00", x"00", x"49", x"75", x"5A", x"76", x"79", x"3D", x"3D", x"3D", x"5D", x"76", x"24", x"00", x"00", x"00", x"00", x"00", x"48", x"71", x"5A", x"3D", x"3D", x"3D", x"5D", x"76", x"00", x"00", x"00", x"00", x"24", x"4D", x"7A", x"4D", x"00", x"00", x"49", x"7A", x"3D", x"76", x"00", x"00"),
( x"00", x"00", x"00", x"6D", x"3D", x"39", x"59", x"71", x"71", x"39", x"39", x"6D", x"00", x"00", x"00", x"00", x"7A", x"19", x"5A", x"24", x"24", x"79", x"39", x"59", x"48", x"00", x"00", x"00", x"6D", x"39", x"39", x"71", x"00", x"00", x"00", x"00", x"20", x"7A", x"39", x"39", x"55", x"6D", x"75", x"59", x"76", x"24", x"00", x"00", x"00", x"71", x"39", x"3D", x"6D", x"49", x"75", x"3D", x"39", x"59", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"72", x"39", x"3D", x"19", x"39", x"75", x"71", x"39", x"39", x"39", x"76", x"00", x"00", x"00", x"00", x"00", x"71", x"39", x"59", x"6D", x"71", x"39", x"5D", x"49", x"00", x"00", x"00", x"28", x"7A", x"5A", x"59", x"59", x"39", x"39", x"75", x"4D", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"5A", x"39", x"39", x"55", x"6D", x"75", x"59", x"76", x"00", x"00", x"00", x"00", x"6D", x"39", x"39", x"4D", x"00", x"00", x"49", x"3D", x"19", x"71", x"00", x"00"),
( x"00", x"00", x"24", x"71", x"39", x"18", x"51", x"24", x"71", x"39", x"39", x"6D", x"00", x"00", x"00", x"20", x"7A", x"18", x"7A", x"24", x"24", x"5A", x"19", x"59", x"28", x"00", x"00", x"00", x"6D", x"39", x"39", x"71", x"00", x"00", x"00", x"00", x"28", x"79", x"18", x"59", x"49", x"00", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"6D", x"39", x"39", x"6D", x"71", x"19", x"39", x"55", x"4D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"71", x"39", x"39", x"55", x"39", x"19", x"39", x"55", x"59", x"19", x"71", x"00", x"00", x"00", x"00", x"4D", x"55", x"39", x"6D", x"00", x"71", x"19", x"59", x"49", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"71", x"39", x"19", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"59", x"18", x"59", x"49", x"00", x"24", x"44", x"24", x"00", x"00", x"00", x"00", x"71", x"39", x"39", x"6D", x"24", x"24", x"6D", x"59", x"39", x"71", x"00", x"00"),
( x"00", x"00", x"71", x"35", x"39", x"55", x"6D", x"00", x"6D", x"39", x"39", x"4D", x"00", x"00", x"00", x"24", x"76", x"14", x"75", x"24", x"24", x"75", x"18", x"55", x"28", x"00", x"00", x"00", x"6D", x"39", x"39", x"71", x"00", x"00", x"00", x"49", x"76", x"39", x"35", x"76", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"39", x"39", x"55", x"35", x"15", x"35", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"71", x"19", x"55", x"49", x"76", x"39", x"76", x"6D", x"55", x"14", x"75", x"00", x"00", x"00", x"00", x"75", x"19", x"39", x"71", x"4D", x"71", x"18", x"59", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"39", x"35", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"76", x"35", x"35", x"76", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"39", x"39", x"55", x"56", x"56", x"55", x"39", x"19", x"71", x"00", x"00"),
( x"00", x"00", x"72", x"14", x"55", x"6D", x"24", x"04", x"71", x"35", x"35", x"4D", x"00", x"00", x"00", x"24", x"76", x"14", x"75", x"24", x"24", x"55", x"14", x"55", x"48", x"00", x"00", x"00", x"6D", x"35", x"35", x"71", x"00", x"00", x"00", x"49", x"35", x"14", x"75", x"24", x"00", x"24", x"6D", x"51", x"6D", x"20", x"00", x"00", x"00", x"6D", x"35", x"35", x"55", x"55", x"35", x"35", x"71", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"71", x"15", x"55", x"49", x"24", x"49", x"24", x"49", x"55", x"14", x"71", x"00", x"00", x"00", x"00", x"71", x"35", x"35", x"35", x"35", x"35", x"35", x"55", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"35", x"14", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"35", x"14", x"75", x"24", x"00", x"24", x"71", x"51", x"71", x"00", x"00", x"00", x"00", x"6D", x"35", x"35", x"55", x"55", x"55", x"55", x"35", x"35", x"71", x"00", x"00"),
( x"00", x"00", x"71", x"11", x"35", x"6D", x"49", x"71", x"55", x"35", x"55", x"4D", x"00", x"00", x"00", x"24", x"76", x"10", x"55", x"49", x"49", x"55", x"10", x"55", x"48", x"00", x"00", x"00", x"6D", x"35", x"35", x"71", x"00", x"00", x"00", x"49", x"35", x"10", x"51", x"44", x"49", x"51", x"35", x"15", x"55", x"24", x"00", x"00", x"00", x"6D", x"35", x"35", x"6D", x"49", x"51", x"35", x"35", x"55", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"71", x"15", x"35", x"49", x"00", x"00", x"00", x"49", x"55", x"10", x"72", x"00", x"00", x"00", x"00", x"71", x"15", x"35", x"51", x"6D", x"51", x"14", x"55", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"35", x"15", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"35", x"10", x"51", x"28", x"4D", x"55", x"35", x"11", x"76", x"00", x"00", x"00", x"00", x"6D", x"15", x"35", x"4D", x"24", x"24", x"4D", x"35", x"15", x"71", x"00", x"00"),
( x"00", x"00", x"6D", x"55", x"11", x"31", x"31", x"11", x"10", x"11", x"51", x"49", x"00", x"00", x"00", x"00", x"76", x"31", x"31", x"31", x"35", x"11", x"31", x"72", x"24", x"00", x"00", x"00", x"6D", x"31", x"11", x"71", x"00", x"00", x"00", x"24", x"76", x"31", x"11", x"55", x"31", x"11", x"35", x"71", x"49", x"00", x"00", x"00", x"00", x"6D", x"11", x"31", x"6D", x"00", x"24", x"6D", x"35", x"11", x"51", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"71", x"11", x"31", x"49", x"00", x"00", x"00", x"49", x"35", x"10", x"72", x"00", x"00", x"00", x"00", x"71", x"11", x"31", x"6D", x"00", x"72", x"11", x"35", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"11", x"11", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"28", x"71", x"31", x"31", x"35", x"31", x"11", x"55", x"71", x"49", x"00", x"00", x"00", x"00", x"6D", x"11", x"11", x"6D", x"00", x"00", x"49", x"35", x"11", x"72", x"00", x"00"),
( x"00", x"00", x"00", x"4D", x"72", x"71", x"72", x"71", x"71", x"31", x"51", x"4D", x"00", x"00", x"00", x"00", x"24", x"6D", x"71", x"71", x"71", x"71", x"6D", x"24", x"00", x"00", x"00", x"00", x"49", x"72", x"72", x"4D", x"00", x"00", x"00", x"00", x"24", x"71", x"72", x"71", x"71", x"71", x"4D", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"72", x"71", x"49", x"00", x"00", x"24", x"71", x"72", x"4D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"71", x"71", x"24", x"00", x"00", x"00", x"24", x"72", x"71", x"6D", x"00", x"00", x"00", x"00", x"4D", x"72", x"71", x"28", x"00", x"6D", x"72", x"72", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"71", x"71", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"71", x"71", x"72", x"71", x"72", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"72", x"71", x"49", x"00", x"00", x"48", x"72", x"72", x"6D", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"00", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"20", x"04", x"20", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"71", x"7A", x"7A", x"7A", x"71", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"76", x"7A", x"7A", x"7A", x"6D", x"00", x"00", x"00", x"00", x"00", x"04", x"4D", x"7A", x"71", x"49", x"00", x"00", x"49", x"71", x"76", x"24", x"00", x"00", x"00", x"00", x"00", x"48", x"49", x"24", x"6D", x"7A", x"7A", x"7A", x"7A", x"76", x"24", x"00", x"00", x"00", x"00", x"00", x"24", x"71", x"7A", x"7A", x"7A", x"71", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"71", x"7A", x"7A", x"7A", x"76", x"24", x"00", x"00", x"00", x"00", x"00", x"4D", x"7A", x"4D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"4D", x"76", x"7A", x"7A", x"7A", x"4D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"7A", x"3D", x"3D", x"59", x"3D", x"3D", x"7A", x"24", x"00", x"00", x"00", x"00", x"4D", x"76", x"59", x"3D", x"5D", x"59", x"3D", x"5A", x"4D", x"00", x"00", x"00", x"00", x"4D", x"5D", x"3D", x"1D", x"7A", x"20", x"24", x"7A", x"39", x"5A", x"24", x"00", x"00", x"00", x"4D", x"76", x"5E", x"5D", x"59", x"59", x"3D", x"59", x"59", x"5A", x"4D", x"00", x"00", x"00", x"00", x"24", x"71", x"7A", x"3D", x"3D", x"59", x"3D", x"3D", x"76", x"00", x"00", x"00", x"00", x"00", x"24", x"71", x"79", x"3D", x"3D", x"59", x"3D", x"3D", x"76", x"00", x"00", x"00", x"00", x"6D", x"5D", x"3D", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"76", x"5D", x"3D", x"3D", x"59", x"59", x"5D", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"59", x"19", x"59", x"71", x"49", x"71", x"75", x"71", x"24", x"00", x"00", x"00", x"00", x"76", x"19", x"39", x"55", x"49", x"71", x"39", x"39", x"4D", x"00", x"00", x"00", x"00", x"71", x"39", x"39", x"38", x"59", x"71", x"4D", x"59", x"19", x"55", x"24", x"00", x"00", x"00", x"71", x"76", x"55", x"75", x"59", x"18", x"59", x"49", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"4D", x"39", x"39", x"59", x"51", x"49", x"59", x"19", x"75", x"04", x"00", x"00", x"00", x"00", x"49", x"59", x"19", x"59", x"71", x"49", x"59", x"18", x"7A", x"24", x"00", x"00", x"00", x"6D", x"39", x"39", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"76", x"39", x"39", x"75", x"4D", x"24", x"49", x"76", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"59", x"14", x"55", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"45", x"76", x"18", x"39", x"4D", x"00", x"71", x"18", x"39", x"6D", x"00", x"00", x"00", x"00", x"6D", x"39", x"38", x"38", x"18", x"59", x"6D", x"55", x"19", x"55", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"75", x"18", x"59", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"59", x"18", x"71", x"24", x"4D", x"59", x"14", x"55", x"24", x"00", x"00", x"00", x"00", x"6D", x"39", x"18", x"55", x"24", x"24", x"59", x"18", x"75", x"24", x"00", x"00", x"00", x"51", x"39", x"39", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"76", x"18", x"39", x"71", x"49", x"28", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"59", x"35", x"55", x"72", x"00", x"00", x"20", x"24", x"00", x"00", x"00", x"00", x"00", x"71", x"35", x"35", x"55", x"49", x"00", x"71", x"15", x"35", x"6D", x"00", x"00", x"00", x"00", x"4D", x"39", x"34", x"55", x"55", x"35", x"71", x"55", x"14", x"55", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"75", x"14", x"55", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"39", x"14", x"75", x"71", x"35", x"35", x"35", x"71", x"00", x"00", x"00", x"00", x"49", x"55", x"35", x"55", x"71", x"00", x"24", x"55", x"14", x"76", x"24", x"00", x"00", x"00", x"6D", x"35", x"35", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"55", x"35", x"35", x"35", x"56", x"72", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"35", x"15", x"71", x"00", x"04", x"49", x"71", x"55", x"71", x"24", x"00", x"00", x"00", x"51", x"14", x"51", x"49", x"20", x"24", x"71", x"14", x"35", x"6D", x"00", x"00", x"00", x"00", x"4D", x"35", x"14", x"6D", x"6D", x"15", x"14", x"34", x"34", x"55", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"75", x"14", x"55", x"48", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"35", x"34", x"35", x"35", x"14", x"51", x"6D", x"24", x"00", x"00", x"00", x"00", x"49", x"35", x"35", x"71", x"04", x"24", x"49", x"55", x"14", x"75", x"24", x"00", x"00", x"00", x"6D", x"35", x"15", x"71", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"6D", x"71", x"51", x"55", x"15", x"35", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"31", x"11", x"51", x"4D", x"6D", x"51", x"11", x"11", x"51", x"24", x"00", x"00", x"00", x"71", x"10", x"51", x"4D", x"4D", x"51", x"31", x"11", x"55", x"49", x"00", x"00", x"00", x"00", x"6D", x"31", x"11", x"6D", x"24", x"71", x"31", x"10", x"10", x"51", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"75", x"10", x"55", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"35", x"10", x"51", x"71", x"10", x"31", x"51", x"49", x"00", x"00", x"00", x"00", x"49", x"35", x"11", x"51", x"4D", x"51", x"35", x"11", x"31", x"72", x"24", x"00", x"00", x"00", x"6D", x"31", x"10", x"51", x"4D", x"4D", x"4D", x"6D", x"49", x"00", x"00", x"00", x"24", x"55", x"31", x"51", x"6D", x"51", x"11", x"31", x"55", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"28", x"71", x"31", x"31", x"31", x"31", x"31", x"51", x"6D", x"24", x"00", x"00", x"00", x"00", x"4D", x"56", x"31", x"31", x"31", x"11", x"51", x"72", x"4D", x"00", x"00", x"00", x"00", x"00", x"6D", x"31", x"11", x"71", x"00", x"28", x"71", x"31", x"11", x"51", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"76", x"11", x"51", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"31", x"11", x"71", x"49", x"72", x"31", x"11", x"72", x"00", x"00", x"00", x"00", x"24", x"72", x"31", x"31", x"31", x"31", x"31", x"55", x"71", x"24", x"00", x"00", x"00", x"00", x"51", x"31", x"31", x"31", x"31", x"31", x"31", x"76", x"4D", x"00", x"00", x"00", x"24", x"71", x"31", x"31", x"31", x"11", x"55", x"71", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"6D", x"6D", x"6D", x"6D", x"44", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6D", x"6D", x"6D", x"6D", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"6D", x"49", x"00", x"00", x"24", x"6D", x"6D", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"6D", x"4D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"6D", x"49", x"00", x"24", x"4D", x"6D", x"49", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"6D", x"6D", x"6D", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6D", x"6D", x"6D", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);

constant SELECTOR_X_size : integer := 16;
constant SELECTOR_Y_size : integer := 16;
type SELECTOR_color_array is array(0 to SELECTOR_Y_size - 1 , 0 to SELECTOR_X_size - 1) of std_logic_vector(7 downto 0);
type SELECTOR_bmp_array is array(0 to SELECTOR_Y_size - 1 , 0 to SELECTOR_X_size - 1) of std_logic;
constant SELECTOR_colors: SELECTOR_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"4D", x"51", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"04", x"49", x"5A", x"7E", x"51", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"04", x"4D", x"5A", x"5E", x"5E", x"5E", x"51", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"24", x"49", x"5A", x"5E", x"59", x"59", x"59", x"5A", x"51", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"4D", x"5A", x"59", x"39", x"39", x"39", x"39", x"39", x"5A", x"51", x"24", x"00", x"00"),
( x"00", x"00", x"49", x"56", x"5A", x"39", x"39", x"38", x"38", x"38", x"39", x"59", x"5A", x"51", x"24", x"00"),
( x"00", x"49", x"56", x"5A", x"39", x"39", x"38", x"38", x"34", x"34", x"38", x"59", x"5A", x"5A", x"4D", x"00"),
( x"00", x"28", x"56", x"5A", x"55", x"35", x"34", x"34", x"34", x"34", x"34", x"35", x"5A", x"56", x"4D", x"00"),
( x"00", x"00", x"28", x"56", x"56", x"35", x"35", x"34", x"34", x"34", x"35", x"35", x"56", x"4D", x"04", x"00"),
( x"00", x"00", x"00", x"49", x"56", x"55", x"35", x"35", x"35", x"35", x"35", x"56", x"4D", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"49", x"52", x"36", x"35", x"35", x"35", x"56", x"4D", x"24", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"20", x"29", x"56", x"56", x"56", x"56", x"4D", x"24", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"20", x"29", x"52", x"56", x"4D", x"24", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"29", x"4D", x"24", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"));

constant CONTROLS_MOVEMENT_KEYS2_X_size : integer := 78;
constant CONTROLS_MOVEMENT_KEYS2_Y_size : integer := 32;
type CONTROLS_MOVEMENT_KEYS2_color_array is array(0 to CONTROLS_MOVEMENT_KEYS2_Y_size - 1 , 0 to CONTROLS_MOVEMENT_KEYS2_X_size - 1) of std_logic_vector(7 downto 0);
constant CONTROLS_MOVEMENT_KEYS2_colors: CONTROLS_MOVEMENT_KEYS2_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"DB", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"B6", x"DB", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"DB", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"00"),
( x"00", x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24"),
( x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92"),
( x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB"),
( x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB"),
( x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB"),
( x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB"),
( x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"6D", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB"),
( x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB"),
( x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB"),
( x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB"),
( x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB"),
( x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92"),
( x"00", x"49", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"B6", x"24"),
( x"00", x"00", x"24", x"49", x"24", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"24", x"24", x"24", x"24", x"24", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"49", x"24", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"24", x"24", x"24", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"49", x"24", x"00")
);


constant CONTROLS_KICK_X_size : integer := 47;
constant CONTROLS_KICK_Y_size : integer := 9;
type CONTROLS_KICK_color_array is array(0 to CONTROLS_KICK_Y_size - 1 , 0 to CONTROLS_KICK_X_size - 1) of std_logic_vector(7 downto 0);
constant CONTROLS_KICK_colors: CONTROLS_KICK_color_array := (
( x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"00"),
( x"00", x"08", x"0C", x"0C", x"00", x"00", x"00", x"04", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"0C", x"0C", x"08", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"04", x"00", x"00", x"04", x"08", x"0C", x"08", x"00"),
( x"00", x"08", x"0C", x"08", x"00", x"04", x"08", x"0C", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"08", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"00", x"00", x"08", x"0C", x"0C", x"04", x"00", x"00"),
( x"00", x"08", x"0C", x"08", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"08", x"04", x"04", x"0C", x"0C", x"00", x"00", x"00", x"00"),
( x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"00"),
( x"00", x"04", x"08", x"08", x"00", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"04", x"08", x"08", x"08", x"00", x"00", x"00"),
( x"00", x"04", x"08", x"04", x"00", x"00", x"04", x"04", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"04", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"04", x"08", x"08", x"04", x"00"),
( x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"04", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);


constant CONTROLS_PUNCH_X_size : integer := 70;
constant CONTROLS_PUNCH_Y_size : integer := 9;
type CONTROLS_PUNCH_color_array is array(0 to CONTROLS_PUNCH_Y_size - 1 , 0 to CONTROLS_PUNCH_X_size - 1) of std_logic_vector(7 downto 0);
constant CONTROLS_PUNCH_colors: CONTROLS_PUNCH_color_array := (
( x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"04"),
( x"00", x"00", x"08", x"0C", x"10", x"0C", x"0C", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"04", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0C", x"08", x"00", x"00", x"00", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"0C", x"0C", x"08", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"04"),
( x"08", x"08", x"0C", x"0C", x"04", x"00", x"04", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"30", x"04", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"0C", x"0C", x"04", x"00", x"00", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"08", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0C", x"00", x"00", x"00", x"00", x"08", x"10", x"08", x"04"),
( x"08", x"0C", x"0C", x"04", x"00", x"00", x"04", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"04", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"08", x"0C", x"0C", x"0C", x"00", x"00", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"04"),
( x"04", x"08", x"0C", x"04", x"00", x"04", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"0C", x"04", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"08", x"08", x"0C", x"00", x"00", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"08", x"08", x"08", x"04", x"08", x"0C", x"08", x"04"),
( x"04", x"08", x"08", x"08", x"08", x"0C", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"08", x"08", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"04"),
( x"04", x"08", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"04", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"04", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"04"),
( x"04", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"04", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"00", x"04", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"04", x"00", x"04", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"04"),
( x"04", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00")
);



constant CONTROLS_MOVEMENT_X_size : integer := 100;
constant CONTROLS_MOVEMENT_Y_size : integer := 8;
type CONTROLS_MOVEMENT_color_array is array(0 to CONTROLS_MOVEMENT_Y_size - 1 , 0 to CONTROLS_MOVEMENT_X_size - 1) of std_logic_vector(7 downto 0);
constant CONTROLS_MOVEMENT_colors: CONTROLS_MOVEMENT_color_array := (
( x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"04"),
( x"04", x"0C", x"10", x"08", x"00", x"00", x"00", x"04", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"0C", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"08", x"10", x"08", x"00", x"00", x"00", x"08", x"10", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"0C", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"10", x"0C", x"04", x"00", x"00", x"04", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"10", x"0C", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"08", x"00", x"00", x"08", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"08", x"0C", x"0C", x"08", x"04", x"00"),
( x"08", x"0C", x"0C", x"0C", x"0C", x"04", x"08", x"2C", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"30", x"0C", x"04", x"00", x"08", x"30", x"04", x"00", x"00", x"00", x"00", x"08", x"10", x"04", x"00", x"00", x"00", x"0C", x"10", x"00", x"00", x"00", x"00", x"00", x"08", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"2C", x"0C", x"0C", x"0C", x"08", x"04", x"0C", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"0C", x"04", x"00", x"08", x"30", x"04", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"0C", x"0C", x"00", x"00", x"00", x"00"),
( x"04", x"0C", x"08", x"00", x"0C", x"30", x"04", x"04", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"08", x"10", x"08", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"08", x"10", x"04", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"08", x"04", x"08", x"10", x"08", x"04", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"0C", x"0C", x"00", x"04", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00", x"00", x"00", x"00"),
( x"04", x"0C", x"04", x"00", x"04", x"04", x"00", x"00", x"0C", x"08", x"00", x"00", x"00", x"00", x"04", x"0C", x"08", x"04", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"04", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"08", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00", x"00", x"04", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0C", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"08", x"04", x"08", x"04", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"00", x"00", x"00", x"00"),
( x"04", x"0C", x"04", x"00", x"00", x"00", x"00", x"04", x"0C", x"08", x"00", x"00", x"00", x"00", x"04", x"0C", x"04", x"00", x"00", x"00", x"04", x"0C", x"04", x"00", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"08", x"0C", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00"),
( x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"04", x"0C", x"08", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"04", x"04", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"04", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00"),
( x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00")
);

constant CONTROLS_ATTACKS_KEYS_X_size : integer := 18;
constant CONTROLS_ATTACKS_KEYS_Y_size : integer := 70;
type CONTROLS_ATTACKS_KEYS_color_array is array(0 to CONTROLS_ATTACKS_KEYS_Y_size - 1 , 0 to CONTROLS_ATTACKS_KEYS_X_size - 1) of std_logic_vector(7 downto 0);
constant CONTROLS_ATTACKS_KEYS_colors: CONTROLS_ATTACKS_KEYS_color_array := (
( x"00", x"49", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"00", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00"),
( x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"6D", x"6D", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"DB", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00"),
( x"24", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"B6", x"24", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"00", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"DB", x"B6", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"92", x"6D", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24"),
( x"00", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"92", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"49", x"92", x"B6", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"B6", x"B6", x"6D", x"00"),
( x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"6D", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"49", x"6D", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"49", x"6D", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"6D", x"92", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"6D", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49"),
( x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"49", x"00")
);

constant CONTROLS_ATTACKS_KEYS2_X_size : integer := 22;
constant CONTROLS_ATTACKS_KEYS2_Y_size : integer := 80;
type CONTROLS_ATTACKS_KEYS2_color_array is array(0 to CONTROLS_ATTACKS_KEYS2_Y_size - 1 , 0 to CONTROLS_ATTACKS_KEYS2_X_size - 1) of std_logic_vector(7 downto 0);
constant CONTROLS_ATTACKS_KEYS2_colors: CONTROLS_ATTACKS_KEYS2_color_array := (
( x"00", x"24", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"49", x"00", x"00", x"00"),
( x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"92", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"92", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00"),
( x"00", x"24", x"49", x"6D", x"49", x"6D", x"49", x"6D", x"49", x"6D", x"6D", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"6D", x"24", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"00", x"00"),
( x"00", x"6D", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"6D", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"6D", x"92", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00"),
( x"00", x"00", x"49", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"49", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"00", x"00"),
( x"00", x"00", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24"),
( x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"49", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"92", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"00", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"00", x"00", x"00", x"49", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"49", x"00")
);

constant CONTROLS_SHOOT_X_size : integer := 70;
constant CONTROLS_SHOOT_Y_size : integer := 9;
type CONTROLS_SHOOT_color_array is array(0 to CONTROLS_SHOOT_Y_size - 1 , 0 to CONTROLS_SHOOT_X_size - 1) of std_logic_vector(7 downto 0);
constant CONTROLS_SHOOT_colors: CONTROLS_SHOOT_color_array := (
( x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"08", x"04"),
( x"00", x"00", x"00", x"08", x"0C", x"0C", x"08", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"08", x"0C", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0C", x"0C", x"0C", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"08", x"0C", x"0C", x"08", x"0C", x"04", x"00"),
( x"00", x"04", x"0C", x"0C", x"08", x"00", x"00", x"00", x"04", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0C", x"00", x"00", x"00", x"00", x"0C", x"10", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"0C", x"04", x"00", x"04", x"10", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"0C", x"08", x"00", x"00", x"08", x"10", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"04", x"08", x"08", x"0C", x"0C", x"08", x"00", x"00", x"00", x"00"),
( x"00", x"04", x"0C", x"0C", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"0C", x"0C", x"08", x"00", x"00", x"04", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"10", x"0C", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00"),
( x"00", x"04", x"0C", x"0C", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"04", x"08", x"08", x"08", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"0C", x"04", x"00", x"00", x"04", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"00", x"00", x"04", x"0C", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"0C", x"08", x"00", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"0C", x"08", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"08", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"00", x"00", x"00", x"00", x"08", x"0C", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00"),
( x"08", x"08", x"08", x"04", x"04", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"08", x"08", x"04", x"04", x"04", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"04", x"04", x"04", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00"),
( x"00", x"04", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"08", x"08", x"08", x"04", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"04", x"08", x"04", x"00", x"00", x"00", x"00")
);


constant CONTROLS_MOVEMENT_KEYS_X_size : integer := 67;
constant CONTROLS_MOVEMENT_KEYS_Y_size : integer := 43;
type CONTROLS_MOVEMENT_KEYS_color_array is array(0 to CONTROLS_MOVEMENT_KEYS_Y_size - 1 , 0 to CONTROLS_MOVEMENT_KEYS_X_size - 1) of std_logic_vector(7 downto 0);

constant CONTROLS_MOVEMENT_KEYS_colors: CONTROLS_MOVEMENT_KEYS_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"FF", x"92", x"B6", x"DB", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"DB", x"49", x"6D", x"B6", x"49", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"6D", x"6D", x"6D", x"6D", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"20", x"92", x"6D", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"DB", x"92", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"DB", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00"),
( x"24", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"92", x"24", x"00", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"49", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"49", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"92", x"B6", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"6D", x"B6", x"49", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"92", x"92", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"24", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"92", x"FF", x"92", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"69", x"49", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"92", x"FF", x"6D", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"92", x"8E", x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"6D", x"49", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"49", x"6D", x"49", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"FF", x"FF", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"92", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"92", x"92", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"49", x"00"),
( x"6D", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"24", x"00"),
( x"24", x"B6", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"DB", x"49", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6", x"00", x"00"),
( x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"00", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00")
);


constant CONTROLS_PLAYER2_X_size : integer := 70;
constant CONTROLS_PLAYER2_Y_size : integer := 9;
type CONTROLS_PLAYER2_color_array is array(0 to CONTROLS_PLAYER2_Y_size - 1 , 0 to CONTROLS_PLAYER2_X_size - 1) of std_logic_vector(7 downto 0);

constant CONTROLS_PLAYER2_colors: CONTROLS_PLAYER2_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"DB", x"DB", x"DB", x"B6", x"49", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"FF", x"DB", x"B6", x"B6", x"FF", x"FF", x"92", x"00"),
( x"00", x"00", x"49", x"92", x"6D", x"00", x"00", x"00", x"00", x"00", x"49", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"24", x"00", x"00", x"00", x"24", x"49", x"00", x"00", x"00", x"49", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"6D", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"49", x"00", x"00", x"00", x"B6", x"FF", x"B6", x"00"),
( x"24", x"B6", x"FF", x"DB", x"FF", x"B6", x"00", x"00", x"00", x"49", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"DB", x"FF", x"FF", x"24", x"00", x"00", x"6D", x"FF", x"49", x"00", x"B6", x"FF", x"24", x"00", x"00", x"00", x"92", x"FF", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"92", x"FF", x"DB", x"DB", x"FF", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"B6", x"00"),
( x"92", x"FF", x"49", x"00", x"FF", x"DB", x"00", x"00", x"00", x"6D", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"B6", x"00", x"92", x"FF", x"24", x"00", x"00", x"49", x"DB", x"FF", x"DB", x"FF", x"B6", x"00", x"00", x"00", x"49", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"92", x"00", x"92", x"FF", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"24", x"00"),
( x"6D", x"FF", x"92", x"B6", x"FF", x"92", x"00", x"00", x"00", x"6D", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"B6", x"24", x"DB", x"FF", x"24", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"DB", x"00", x"00", x"00", x"00", x"49", x"FF", x"DB", x"B6", x"92", x"00", x"00", x"00", x"00", x"6D", x"FF", x"92", x"92", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"B6", x"24", x"00", x"00"),
( x"6D", x"FF", x"DB", x"DB", x"49", x"00", x"00", x"00", x"00", x"6D", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"DB", x"B6", x"FF", x"FF", x"24", x"00", x"00", x"00", x"00", x"DB", x"FF", x"24", x"00", x"00", x"00", x"00", x"49", x"FF", x"B6", x"24", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"DB", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"92", x"49", x"24", x"49", x"24"),
( x"92", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"DB", x"DB", x"92", x"00", x"00", x"00", x"49", x"FF", x"92", x"00", x"B6", x"FF", x"49", x"00", x"00", x"00", x"00", x"B6", x"FF", x"49", x"00", x"00", x"00", x"00", x"49", x"FF", x"DB", x"B6", x"DB", x"92", x"00", x"00", x"00", x"6D", x"FF", x"6D", x"6D", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"FF", x"6D"),
( x"24", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"6D", x"6D", x"00", x"00", x"00", x"00", x"00", x"6D", x"24", x"00", x"24", x"49", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6D", x"6D", x"6D", x"24", x"00", x"00", x"00", x"00", x"49", x"24", x"00", x"24", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"49", x"49", x"49", x"49", x"49", x"49", x"24", x"00")
);


constant CONTROLS_PLAYER1_X_size : integer := 70;
constant CONTROLS_PLAYER1_Y_size : integer := 9;
type CONTROLS_PLAYER1_color_array is array(0 to CONTROLS_PLAYER1_Y_size - 1 , 0 to CONTROLS_PLAYER1_X_size - 1) of std_logic_vector(7 downto 0);

constant CONTROLS_PLAYER1_colors: CONTROLS_PLAYER1_color_array := (
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"B6", x"DB", x"B6", x"00", x"00"),
( x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"DB", x"00", x"00"),
( x"00", x"00", x"24", x"92", x"6D", x"24", x"00", x"00", x"00", x"00", x"24", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"49", x"00", x"00", x"00", x"00", x"49", x"24", x"00", x"00", x"00", x"49", x"00", x"00", x"00", x"00", x"00", x"49", x"92", x"92", x"49", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"49", x"49", x"DB", x"FF", x"DB", x"00", x"00"),
( x"24", x"B6", x"FF", x"DB", x"FF", x"FF", x"24", x"00", x"00", x"00", x"DB", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"DB", x"DB", x"FF", x"92", x"00", x"00", x"00", x"B6", x"FF", x"24", x"00", x"DB", x"FF", x"00", x"00", x"00", x"24", x"B6", x"FF", x"DB", x"B6", x"49", x"00", x"00", x"00", x"00", x"92", x"FF", x"DB", x"DB", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"DB", x"00", x"00"),
( x"49", x"FF", x"92", x"00", x"B6", x"FF", x"24", x"00", x"00", x"00", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"6D", x"DB", x"00", x"00", x"FF", x"B6", x"00", x"00", x"00", x"6D", x"FF", x"FF", x"DB", x"FF", x"B6", x"00", x"00", x"00", x"92", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"B6", x"00", x"6D", x"FF", x"6D", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"DB", x"00", x"00"),
( x"6D", x"FF", x"92", x"6D", x"FF", x"DB", x"00", x"00", x"00", x"00", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"49", x"6D", x"FF", x"92", x"00", x"00", x"00", x"00", x"B6", x"FF", x"FF", x"B6", x"00", x"00", x"00", x"00", x"92", x"FF", x"DB", x"B6", x"6D", x"00", x"00", x"00", x"00", x"49", x"FF", x"B6", x"6D", x"FF", x"DB", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"B6", x"FF", x"DB", x"00", x"00"),
( x"49", x"FF", x"DB", x"DB", x"6D", x"00", x"00", x"00", x"00", x"00", x"FF", x"DB", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"DB", x"DB", x"FF", x"92", x"00", x"00", x"00", x"00", x"24", x"FF", x"FF", x"00", x"00", x"00", x"00", x"00", x"92", x"FF", x"92", x"24", x"00", x"00", x"00", x"00", x"00", x"49", x"FF", x"FF", x"FF", x"FF", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"DB", x"FF", x"DB", x"49", x"24"),
( x"49", x"FF", x"92", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"FF", x"FF", x"DB", x"DB", x"B6", x"49", x"00", x"00", x"00", x"FF", x"FF", x"00", x"24", x"FF", x"B6", x"00", x"00", x"00", x"00", x"00", x"DB", x"FF", x"24", x"00", x"00", x"00", x"00", x"92", x"FF", x"DB", x"B6", x"DB", x"6D", x"00", x"00", x"00", x"49", x"FF", x"92", x"49", x"FF", x"FF", x"49", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"92", x"FF", x"FF", x"FF", x"FF", x"FF", x"B6"),
( x"24", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"49", x"6D", x"6D", x"6D", x"49", x"00", x"00", x"00", x"00", x"49", x"49", x"00", x"00", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"49", x"49", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"6D", x"6D", x"6D", x"24", x"00", x"00", x"00", x"24", x"6D", x"49", x"00", x"24", x"6D", x"24", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"24", x"6D", x"49", x"49", x"49", x"49", x"49", x"49")
);


constant press_Start_X	: integer := 190;
constant press_End_X 	: integer := press_Start_X + press_S_X_size;
constant press_Start_Y 	: integer := 350;
constant press_End_Y 	: integer := press_Start_Y + press_S_Y_size;

constant OPTIONS_Start_X : integer := 250;
constant OPTIONS_End_X : integer := OPTIONS_Start_X + OPTIONS_X_size;

constant OPTIONS_Start_Y : integer :=  320;
constant OPTIONS_End_Y : integer := OPTIONS_Start_Y + OPTIONS_Y_size;

constant CONTROLS_MENU_Start_X : integer := 187;
constant CONTROLS_MENU_End_X: integer := CONTROLS_MENU_Start_X + CONTROLS_MOVEMENT_KEYS_X_size + CONTROLS_MOVEMENT_X_size + 20 + CONTROLS_MOVEMENT_KEYS2_X_size ;

constant CONTROLS_MENU_Start_Y : integer := OPTIONS_Start_Y;
constant CONTROLS_MENU_End_Y : integer := OPTIONS_Start_Y + 140;

constant CONTROLS_MENU_MOVEMENT_KEYS1_Start_X : integer := CONTROLS_MENU_Start_X;
constant CONTROLS_MENU_MOVEMENT_KEYS1_End_X : integer := CONTROLS_MENU_Start_X + CONTROLS_MOVEMENT_KEYS_X_size;

constant CONTROLS_MENU_MOVEMENT_KEYS1_Start_Y : integer := CONTROLS_MENU_Start_Y + CONTROLS_PLAYER1_Y_size + 4;
constant CONTROLS_MENU_MOVEMENT_KEYS1_End_Y : integer := CONTROLS_MENU_MOVEMENT_KEYS1_Start_Y + CONTROLS_MOVEMENT_KEYS_Y_size;

constant CONTROLS_MENU_MOVEMENT_KEYS2_Start_X : integer := CONTROLS_MENU_MOVEMENT_KEYS1_End_X + CONTROLS_MOVEMENT_X_size + 20;
constant CONTROLS_MENU_MOVEMENT_KEYS2_End_X : integer := CONTROLS_MENU_MOVEMENT_KEYS2_Start_X + CONTROLS_MOVEMENT_KEYS2_X_size;

constant CONTROLS_MENU_MOVEMENT_KEYS2_Start_Y : integer := CONTROLS_MENU_Start_Y + CONTROLS_PLAYER2_Y_size + 4;
constant CONTROLS_MENU_MOVEMENT_KEYS2_End_Y : integer := CONTROLS_MENU_MOVEMENT_KEYS2_Start_Y + CONTROLS_MOVEMENT_KEYS2_Y_size;

constant CONTROLS_MENU_ATTACK_KEYS1_Start_X : integer := CONTROLS_MENU_MOVEMENT_KEYS1_Start_X + 20;
constant CONTROLS_MENU_ATTACK_KEYS1_End_X : integer := CONTROLS_MENU_ATTACK_KEYS1_Start_X + CONTROLS_ATTACKS_KEYS_X_size;

constant CONTROLS_MENU_ATTACK_KEYS1_Start_Y : integer := CONTROLS_MENU_MOVEMENT_KEYS1_End_Y + 4;
constant CONTROLS_MENU_ATTACK_KEYS1_End_Y : integer := CONTROLS_MENU_ATTACK_KEYS1_Start_Y + CONTROLS_ATTACKS_KEYS_Y_size;

constant CONTROLS_MENU_ATTACK_KEYS2_Start_X : integer := CONTROLS_MENU_MOVEMENT_KEYS2_Start_X + 30;
constant CONTROLS_MENU_ATTACK_KEYS2_End_X : integer := CONTROLS_MENU_ATTACK_KEYS2_Start_X + CONTROLS_ATTACKS_KEYS2_X_size;

constant CONTROLS_MENU_ATTACK_KEYS2_Start_Y : integer := CONTROLS_MENU_MOVEMENT_KEYS2_End_Y + 10;
constant CONTROLS_MENU_ATTACK_KEYS2_End_Y : integer := CONTROLS_MENU_ATTACK_KEYS2_Start_Y + CONTROLS_ATTACKS_KEYS2_Y_size;

end MAIN_MENU_PCKG;